module PartialProductGenerator(
  output [0:0] pp_0,
  output [1:0] pp_1,
  output [2:0] pp_2,
  output [3:0] pp_3,
  output [4:0] pp_4,
  output [5:0] pp_5,
  output [6:0] pp_6,
  output [7:0] pp_7,
  output [8:0] pp_8,
  output [9:0] pp_9,
  output [10:0] pp_10,
  output [11:0] pp_11,
  output [12:0] pp_12,
  output [13:0] pp_13,
  output [14:0] pp_14,
  output [15:0] pp_15,
  output [14:0] pp_16,
  output [13:0] pp_17,
  output [12:0] pp_18,
  output [11:0] pp_19,
  output [10:0] pp_20,
  output [9:0] pp_21,
  output [8:0] pp_22,
  output [7:0] pp_23,
  output [6:0] pp_24,
  output [5:0] pp_25,
  output [4:0] pp_26,
  output [3:0] pp_27,
  output [2:0] pp_28,
  output [1:0] pp_29,
  output [0:0] pp_30,
  input [15:0] multiplicand,
  input [15:0] multiplier
);
  assign pp_0[0] = multiplicand[0] & multiplier[0];
  assign pp_1[0] = multiplicand[0] & multiplier[1];
  assign pp_1[1] = multiplicand[1] & multiplier[0];
  assign pp_2[0] = multiplicand[0] & multiplier[2];
  assign pp_2[1] = multiplicand[1] & multiplier[1];
  assign pp_2[2] = multiplicand[2] & multiplier[0];
  assign pp_3[0] = multiplicand[0] & multiplier[3];
  assign pp_3[1] = multiplicand[1] & multiplier[2];
  assign pp_3[2] = multiplicand[2] & multiplier[1];
  assign pp_3[3] = multiplicand[3] & multiplier[0];
  assign pp_4[0] = multiplicand[0] & multiplier[4];
  assign pp_4[1] = multiplicand[1] & multiplier[3];
  assign pp_4[2] = multiplicand[2] & multiplier[2];
  assign pp_4[3] = multiplicand[3] & multiplier[1];
  assign pp_4[4] = multiplicand[4] & multiplier[0];
  assign pp_5[0] = multiplicand[0] & multiplier[5];
  assign pp_5[1] = multiplicand[1] & multiplier[4];
  assign pp_5[2] = multiplicand[2] & multiplier[3];
  assign pp_5[3] = multiplicand[3] & multiplier[2];
  assign pp_5[4] = multiplicand[4] & multiplier[1];
  assign pp_5[5] = multiplicand[5] & multiplier[0];
  assign pp_6[0] = multiplicand[0] & multiplier[6];
  assign pp_6[1] = multiplicand[1] & multiplier[5];
  assign pp_6[2] = multiplicand[2] & multiplier[4];
  assign pp_6[3] = multiplicand[3] & multiplier[3];
  assign pp_6[4] = multiplicand[4] & multiplier[2];
  assign pp_6[5] = multiplicand[5] & multiplier[1];
  assign pp_6[6] = multiplicand[6] & multiplier[0];
  assign pp_7[0] = multiplicand[0] & multiplier[7];
  assign pp_7[1] = multiplicand[1] & multiplier[6];
  assign pp_7[2] = multiplicand[2] & multiplier[5];
  assign pp_7[3] = multiplicand[3] & multiplier[4];
  assign pp_7[4] = multiplicand[4] & multiplier[3];
  assign pp_7[5] = multiplicand[5] & multiplier[2];
  assign pp_7[6] = multiplicand[6] & multiplier[1];
  assign pp_7[7] = multiplicand[7] & multiplier[0];
  assign pp_8[0] = multiplicand[0] & multiplier[8];
  assign pp_8[1] = multiplicand[1] & multiplier[7];
  assign pp_8[2] = multiplicand[2] & multiplier[6];
  assign pp_8[3] = multiplicand[3] & multiplier[5];
  assign pp_8[4] = multiplicand[4] & multiplier[4];
  assign pp_8[5] = multiplicand[5] & multiplier[3];
  assign pp_8[6] = multiplicand[6] & multiplier[2];
  assign pp_8[7] = multiplicand[7] & multiplier[1];
  assign pp_8[8] = multiplicand[8] & multiplier[0];
  assign pp_9[0] = multiplicand[0] & multiplier[9];
  assign pp_9[1] = multiplicand[1] & multiplier[8];
  assign pp_9[2] = multiplicand[2] & multiplier[7];
  assign pp_9[3] = multiplicand[3] & multiplier[6];
  assign pp_9[4] = multiplicand[4] & multiplier[5];
  assign pp_9[5] = multiplicand[5] & multiplier[4];
  assign pp_9[6] = multiplicand[6] & multiplier[3];
  assign pp_9[7] = multiplicand[7] & multiplier[2];
  assign pp_9[8] = multiplicand[8] & multiplier[1];
  assign pp_9[9] = multiplicand[9] & multiplier[0];
  assign pp_10[0] = multiplicand[0] & multiplier[10];
  assign pp_10[1] = multiplicand[1] & multiplier[9];
  assign pp_10[2] = multiplicand[2] & multiplier[8];
  assign pp_10[3] = multiplicand[3] & multiplier[7];
  assign pp_10[4] = multiplicand[4] & multiplier[6];
  assign pp_10[5] = multiplicand[5] & multiplier[5];
  assign pp_10[6] = multiplicand[6] & multiplier[4];
  assign pp_10[7] = multiplicand[7] & multiplier[3];
  assign pp_10[8] = multiplicand[8] & multiplier[2];
  assign pp_10[9] = multiplicand[9] & multiplier[1];
  assign pp_10[10] = multiplicand[10] & multiplier[0];
  assign pp_11[0] = multiplicand[0] & multiplier[11];
  assign pp_11[1] = multiplicand[1] & multiplier[10];
  assign pp_11[2] = multiplicand[2] & multiplier[9];
  assign pp_11[3] = multiplicand[3] & multiplier[8];
  assign pp_11[4] = multiplicand[4] & multiplier[7];
  assign pp_11[5] = multiplicand[5] & multiplier[6];
  assign pp_11[6] = multiplicand[6] & multiplier[5];
  assign pp_11[7] = multiplicand[7] & multiplier[4];
  assign pp_11[8] = multiplicand[8] & multiplier[3];
  assign pp_11[9] = multiplicand[9] & multiplier[2];
  assign pp_11[10] = multiplicand[10] & multiplier[1];
  assign pp_11[11] = multiplicand[11] & multiplier[0];
  assign pp_12[0] = multiplicand[0] & multiplier[12];
  assign pp_12[1] = multiplicand[1] & multiplier[11];
  assign pp_12[2] = multiplicand[2] & multiplier[10];
  assign pp_12[3] = multiplicand[3] & multiplier[9];
  assign pp_12[4] = multiplicand[4] & multiplier[8];
  assign pp_12[5] = multiplicand[5] & multiplier[7];
  assign pp_12[6] = multiplicand[6] & multiplier[6];
  assign pp_12[7] = multiplicand[7] & multiplier[5];
  assign pp_12[8] = multiplicand[8] & multiplier[4];
  assign pp_12[9] = multiplicand[9] & multiplier[3];
  assign pp_12[10] = multiplicand[10] & multiplier[2];
  assign pp_12[11] = multiplicand[11] & multiplier[1];
  assign pp_12[12] = multiplicand[12] & multiplier[0];
  assign pp_13[0] = multiplicand[0] & multiplier[13];
  assign pp_13[1] = multiplicand[1] & multiplier[12];
  assign pp_13[2] = multiplicand[2] & multiplier[11];
  assign pp_13[3] = multiplicand[3] & multiplier[10];
  assign pp_13[4] = multiplicand[4] & multiplier[9];
  assign pp_13[5] = multiplicand[5] & multiplier[8];
  assign pp_13[6] = multiplicand[6] & multiplier[7];
  assign pp_13[7] = multiplicand[7] & multiplier[6];
  assign pp_13[8] = multiplicand[8] & multiplier[5];
  assign pp_13[9] = multiplicand[9] & multiplier[4];
  assign pp_13[10] = multiplicand[10] & multiplier[3];
  assign pp_13[11] = multiplicand[11] & multiplier[2];
  assign pp_13[12] = multiplicand[12] & multiplier[1];
  assign pp_13[13] = multiplicand[13] & multiplier[0];
  assign pp_14[0] = multiplicand[0] & multiplier[14];
  assign pp_14[1] = multiplicand[1] & multiplier[13];
  assign pp_14[2] = multiplicand[2] & multiplier[12];
  assign pp_14[3] = multiplicand[3] & multiplier[11];
  assign pp_14[4] = multiplicand[4] & multiplier[10];
  assign pp_14[5] = multiplicand[5] & multiplier[9];
  assign pp_14[6] = multiplicand[6] & multiplier[8];
  assign pp_14[7] = multiplicand[7] & multiplier[7];
  assign pp_14[8] = multiplicand[8] & multiplier[6];
  assign pp_14[9] = multiplicand[9] & multiplier[5];
  assign pp_14[10] = multiplicand[10] & multiplier[4];
  assign pp_14[11] = multiplicand[11] & multiplier[3];
  assign pp_14[12] = multiplicand[12] & multiplier[2];
  assign pp_14[13] = multiplicand[13] & multiplier[1];
  assign pp_14[14] = multiplicand[14] & multiplier[0];
  assign pp_15[0] = multiplicand[0] & multiplier[15];
  assign pp_15[1] = multiplicand[1] & multiplier[14];
  assign pp_15[2] = multiplicand[2] & multiplier[13];
  assign pp_15[3] = multiplicand[3] & multiplier[12];
  assign pp_15[4] = multiplicand[4] & multiplier[11];
  assign pp_15[5] = multiplicand[5] & multiplier[10];
  assign pp_15[6] = multiplicand[6] & multiplier[9];
  assign pp_15[7] = multiplicand[7] & multiplier[8];
  assign pp_15[8] = multiplicand[8] & multiplier[7];
  assign pp_15[9] = multiplicand[9] & multiplier[6];
  assign pp_15[10] = multiplicand[10] & multiplier[5];
  assign pp_15[11] = multiplicand[11] & multiplier[4];
  assign pp_15[12] = multiplicand[12] & multiplier[3];
  assign pp_15[13] = multiplicand[13] & multiplier[2];
  assign pp_15[14] = multiplicand[14] & multiplier[1];
  assign pp_15[15] = multiplicand[15] & multiplier[0];
  assign pp_16[0] = multiplicand[1] & multiplier[15];
  assign pp_16[1] = multiplicand[2] & multiplier[14];
  assign pp_16[2] = multiplicand[3] & multiplier[13];
  assign pp_16[3] = multiplicand[4] & multiplier[12];
  assign pp_16[4] = multiplicand[5] & multiplier[11];
  assign pp_16[5] = multiplicand[6] & multiplier[10];
  assign pp_16[6] = multiplicand[7] & multiplier[9];
  assign pp_16[7] = multiplicand[8] & multiplier[8];
  assign pp_16[8] = multiplicand[9] & multiplier[7];
  assign pp_16[9] = multiplicand[10] & multiplier[6];
  assign pp_16[10] = multiplicand[11] & multiplier[5];
  assign pp_16[11] = multiplicand[12] & multiplier[4];
  assign pp_16[12] = multiplicand[13] & multiplier[3];
  assign pp_16[13] = multiplicand[14] & multiplier[2];
  assign pp_16[14] = multiplicand[15] & multiplier[1];
  assign pp_17[0] = multiplicand[2] & multiplier[15];
  assign pp_17[1] = multiplicand[3] & multiplier[14];
  assign pp_17[2] = multiplicand[4] & multiplier[13];
  assign pp_17[3] = multiplicand[5] & multiplier[12];
  assign pp_17[4] = multiplicand[6] & multiplier[11];
  assign pp_17[5] = multiplicand[7] & multiplier[10];
  assign pp_17[6] = multiplicand[8] & multiplier[9];
  assign pp_17[7] = multiplicand[9] & multiplier[8];
  assign pp_17[8] = multiplicand[10] & multiplier[7];
  assign pp_17[9] = multiplicand[11] & multiplier[6];
  assign pp_17[10] = multiplicand[12] & multiplier[5];
  assign pp_17[11] = multiplicand[13] & multiplier[4];
  assign pp_17[12] = multiplicand[14] & multiplier[3];
  assign pp_17[13] = multiplicand[15] & multiplier[2];
  assign pp_18[0] = multiplicand[3] & multiplier[15];
  assign pp_18[1] = multiplicand[4] & multiplier[14];
  assign pp_18[2] = multiplicand[5] & multiplier[13];
  assign pp_18[3] = multiplicand[6] & multiplier[12];
  assign pp_18[4] = multiplicand[7] & multiplier[11];
  assign pp_18[5] = multiplicand[8] & multiplier[10];
  assign pp_18[6] = multiplicand[9] & multiplier[9];
  assign pp_18[7] = multiplicand[10] & multiplier[8];
  assign pp_18[8] = multiplicand[11] & multiplier[7];
  assign pp_18[9] = multiplicand[12] & multiplier[6];
  assign pp_18[10] = multiplicand[13] & multiplier[5];
  assign pp_18[11] = multiplicand[14] & multiplier[4];
  assign pp_18[12] = multiplicand[15] & multiplier[3];
  assign pp_19[0] = multiplicand[4] & multiplier[15];
  assign pp_19[1] = multiplicand[5] & multiplier[14];
  assign pp_19[2] = multiplicand[6] & multiplier[13];
  assign pp_19[3] = multiplicand[7] & multiplier[12];
  assign pp_19[4] = multiplicand[8] & multiplier[11];
  assign pp_19[5] = multiplicand[9] & multiplier[10];
  assign pp_19[6] = multiplicand[10] & multiplier[9];
  assign pp_19[7] = multiplicand[11] & multiplier[8];
  assign pp_19[8] = multiplicand[12] & multiplier[7];
  assign pp_19[9] = multiplicand[13] & multiplier[6];
  assign pp_19[10] = multiplicand[14] & multiplier[5];
  assign pp_19[11] = multiplicand[15] & multiplier[4];
  assign pp_20[0] = multiplicand[5] & multiplier[15];
  assign pp_20[1] = multiplicand[6] & multiplier[14];
  assign pp_20[2] = multiplicand[7] & multiplier[13];
  assign pp_20[3] = multiplicand[8] & multiplier[12];
  assign pp_20[4] = multiplicand[9] & multiplier[11];
  assign pp_20[5] = multiplicand[10] & multiplier[10];
  assign pp_20[6] = multiplicand[11] & multiplier[9];
  assign pp_20[7] = multiplicand[12] & multiplier[8];
  assign pp_20[8] = multiplicand[13] & multiplier[7];
  assign pp_20[9] = multiplicand[14] & multiplier[6];
  assign pp_20[10] = multiplicand[15] & multiplier[5];
  assign pp_21[0] = multiplicand[6] & multiplier[15];
  assign pp_21[1] = multiplicand[7] & multiplier[14];
  assign pp_21[2] = multiplicand[8] & multiplier[13];
  assign pp_21[3] = multiplicand[9] & multiplier[12];
  assign pp_21[4] = multiplicand[10] & multiplier[11];
  assign pp_21[5] = multiplicand[11] & multiplier[10];
  assign pp_21[6] = multiplicand[12] & multiplier[9];
  assign pp_21[7] = multiplicand[13] & multiplier[8];
  assign pp_21[8] = multiplicand[14] & multiplier[7];
  assign pp_21[9] = multiplicand[15] & multiplier[6];
  assign pp_22[0] = multiplicand[7] & multiplier[15];
  assign pp_22[1] = multiplicand[8] & multiplier[14];
  assign pp_22[2] = multiplicand[9] & multiplier[13];
  assign pp_22[3] = multiplicand[10] & multiplier[12];
  assign pp_22[4] = multiplicand[11] & multiplier[11];
  assign pp_22[5] = multiplicand[12] & multiplier[10];
  assign pp_22[6] = multiplicand[13] & multiplier[9];
  assign pp_22[7] = multiplicand[14] & multiplier[8];
  assign pp_22[8] = multiplicand[15] & multiplier[7];
  assign pp_23[0] = multiplicand[8] & multiplier[15];
  assign pp_23[1] = multiplicand[9] & multiplier[14];
  assign pp_23[2] = multiplicand[10] & multiplier[13];
  assign pp_23[3] = multiplicand[11] & multiplier[12];
  assign pp_23[4] = multiplicand[12] & multiplier[11];
  assign pp_23[5] = multiplicand[13] & multiplier[10];
  assign pp_23[6] = multiplicand[14] & multiplier[9];
  assign pp_23[7] = multiplicand[15] & multiplier[8];
  assign pp_24[0] = multiplicand[9] & multiplier[15];
  assign pp_24[1] = multiplicand[10] & multiplier[14];
  assign pp_24[2] = multiplicand[11] & multiplier[13];
  assign pp_24[3] = multiplicand[12] & multiplier[12];
  assign pp_24[4] = multiplicand[13] & multiplier[11];
  assign pp_24[5] = multiplicand[14] & multiplier[10];
  assign pp_24[6] = multiplicand[15] & multiplier[9];
  assign pp_25[0] = multiplicand[10] & multiplier[15];
  assign pp_25[1] = multiplicand[11] & multiplier[14];
  assign pp_25[2] = multiplicand[12] & multiplier[13];
  assign pp_25[3] = multiplicand[13] & multiplier[12];
  assign pp_25[4] = multiplicand[14] & multiplier[11];
  assign pp_25[5] = multiplicand[15] & multiplier[10];
  assign pp_26[0] = multiplicand[11] & multiplier[15];
  assign pp_26[1] = multiplicand[12] & multiplier[14];
  assign pp_26[2] = multiplicand[13] & multiplier[13];
  assign pp_26[3] = multiplicand[14] & multiplier[12];
  assign pp_26[4] = multiplicand[15] & multiplier[11];
  assign pp_27[0] = multiplicand[12] & multiplier[15];
  assign pp_27[1] = multiplicand[13] & multiplier[14];
  assign pp_27[2] = multiplicand[14] & multiplier[13];
  assign pp_27[3] = multiplicand[15] & multiplier[12];
  assign pp_28[0] = multiplicand[13] & multiplier[15];
  assign pp_28[1] = multiplicand[14] & multiplier[14];
  assign pp_28[2] = multiplicand[15] & multiplier[13];
  assign pp_29[0] = multiplicand[14] & multiplier[15];
  assign pp_29[1] = multiplicand[15] & multiplier[14];
  assign pp_30[0] = multiplicand[15] & multiplier[15];
endmodule

`ifndef OP_COMPTREE_FA
`define OP_COMPTREE_FA

module FullAdder(
  input   io_a,
  input   io_b,
  input   io_ci,
  output  io_s,
  output  io_co
);
`ifdef DC
  DW01_add #(1) 
    adder ( .A(io_a), .B(io_b), .CI(io_ci), .SUM(io_s), .CO(io_co) );
`else
  wire  a_xor_b = io_a ^ io_b;
  wire  a_and_b = io_a & io_b;
  wire  a_and_cin = io_a & io_ci;
  wire  b_and_cin = io_b & io_ci;
  wire  _T_1 = a_and_b | b_and_cin;
  assign io_s = a_xor_b ^ io_ci;
  assign io_co = _T_1 | a_and_cin;
`endif
endmodule

`endif


`ifndef OP_COMPTREE_HA
`define OP_COMPTREE_HA

module HalfAdder(
  input   io_a,
  input   io_b,
  output  io_s,
  output  io_co
);
  assign io_s = io_a ^ io_b;
  assign io_co = io_a & io_b;
endmodule

`endif


`ifndef OP_COMPTREE_FT
`define OP_COMPTREE_FT

module FallThrough(
  input  io_a,
  output io_s
);
  assign io_s = io_a;
endmodule

`endif
module CompressorTree(
  input clock,
  input reset,
  input [0:0] io_pp_0,
  input [1:0] io_pp_1,
  input [2:0] io_pp_2,
  input [3:0] io_pp_3,
  input [4:0] io_pp_4,
  input [5:0] io_pp_5,
  input [6:0] io_pp_6,
  input [7:0] io_pp_7,
  input [8:0] io_pp_8,
  input [9:0] io_pp_9,
  input [10:0] io_pp_10,
  input [11:0] io_pp_11,
  input [12:0] io_pp_12,
  input [13:0] io_pp_13,
  input [14:0] io_pp_14,
  input [15:0] io_pp_15,
  input [14:0] io_pp_16,
  input [13:0] io_pp_17,
  input [12:0] io_pp_18,
  input [11:0] io_pp_19,
  input [10:0] io_pp_20,
  input [9:0] io_pp_21,
  input [8:0] io_pp_22,
  input [7:0] io_pp_23,
  input [6:0] io_pp_24,
  input [5:0] io_pp_25,
  input [4:0] io_pp_26,
  input [3:0] io_pp_27,
  input [2:0] io_pp_28,
  input [1:0] io_pp_29,
  input [0:0] io_pp_30,
  output [31:0] io_augend,
  output [31:0] io_addend
);
  wire ft_s0_c0_r0_io_a;
  wire ft_s0_c0_r0_io_s;
  FallThrough ft_s0_c0_r0(
    .io_a(ft_s0_c0_r0_io_a),
    .io_s(ft_s0_c0_r0_io_s)
  );
  wire ft_s1_c0_r0_io_a;
  wire ft_s1_c0_r0_io_s;
  FallThrough ft_s1_c0_r0(
    .io_a(ft_s1_c0_r0_io_a),
    .io_s(ft_s1_c0_r0_io_s)
  );
  wire ft_s2_c0_r0_io_a;
  wire ft_s2_c0_r0_io_s;
  FallThrough ft_s2_c0_r0(
    .io_a(ft_s2_c0_r0_io_a),
    .io_s(ft_s2_c0_r0_io_s)
  );
  wire ft_s3_c0_r0_io_a;
  wire ft_s3_c0_r0_io_s;
  FallThrough ft_s3_c0_r0(
    .io_a(ft_s3_c0_r0_io_a),
    .io_s(ft_s3_c0_r0_io_s)
  );
  wire ft_s4_c0_r0_io_a;
  wire ft_s4_c0_r0_io_s;
  FallThrough ft_s4_c0_r0(
    .io_a(ft_s4_c0_r0_io_a),
    .io_s(ft_s4_c0_r0_io_s)
  );
  wire ft_s5_c0_r0_io_a;
  wire ft_s5_c0_r0_io_s;
  FallThrough ft_s5_c0_r0(
    .io_a(ft_s5_c0_r0_io_a),
    .io_s(ft_s5_c0_r0_io_s)
  );
  wire ft_s6_c0_r0_io_a;
  wire ft_s6_c0_r0_io_s;
  FallThrough ft_s6_c0_r0(
    .io_a(ft_s6_c0_r0_io_a),
    .io_s(ft_s6_c0_r0_io_s)
  );
  wire ft_s7_c0_r0_io_a;
  wire ft_s7_c0_r0_io_s;
  FallThrough ft_s7_c0_r0(
    .io_a(ft_s7_c0_r0_io_a),
    .io_s(ft_s7_c0_r0_io_s)
  );
  wire ft_s8_c0_r0_io_a;
  wire ft_s8_c0_r0_io_s;
  FallThrough ft_s8_c0_r0(
    .io_a(ft_s8_c0_r0_io_a),
    .io_s(ft_s8_c0_r0_io_s)
  );
  wire ha_s0_c1_r0_io_a;
  wire ha_s0_c1_r0_io_b;
  wire ha_s0_c1_r0_io_s;
  wire ha_s0_c1_r0_io_co;
  HalfAdder ha_s0_c1_r0(
    .io_a(ha_s0_c1_r0_io_a),
    .io_b(ha_s0_c1_r0_io_b),
    .io_s(ha_s0_c1_r0_io_s),
    .io_co(ha_s0_c1_r0_io_co)
  );
  wire ft_s1_c1_r0_io_a;
  wire ft_s1_c1_r0_io_s;
  FallThrough ft_s1_c1_r0(
    .io_a(ft_s1_c1_r0_io_a),
    .io_s(ft_s1_c1_r0_io_s)
  );
  wire ft_s2_c1_r0_io_a;
  wire ft_s2_c1_r0_io_s;
  FallThrough ft_s2_c1_r0(
    .io_a(ft_s2_c1_r0_io_a),
    .io_s(ft_s2_c1_r0_io_s)
  );
  wire ft_s3_c1_r0_io_a;
  wire ft_s3_c1_r0_io_s;
  FallThrough ft_s3_c1_r0(
    .io_a(ft_s3_c1_r0_io_a),
    .io_s(ft_s3_c1_r0_io_s)
  );
  wire ft_s4_c1_r0_io_a;
  wire ft_s4_c1_r0_io_s;
  FallThrough ft_s4_c1_r0(
    .io_a(ft_s4_c1_r0_io_a),
    .io_s(ft_s4_c1_r0_io_s)
  );
  wire ft_s5_c1_r0_io_a;
  wire ft_s5_c1_r0_io_s;
  FallThrough ft_s5_c1_r0(
    .io_a(ft_s5_c1_r0_io_a),
    .io_s(ft_s5_c1_r0_io_s)
  );
  wire ft_s6_c1_r0_io_a;
  wire ft_s6_c1_r0_io_s;
  FallThrough ft_s6_c1_r0(
    .io_a(ft_s6_c1_r0_io_a),
    .io_s(ft_s6_c1_r0_io_s)
  );
  wire ft_s7_c1_r0_io_a;
  wire ft_s7_c1_r0_io_s;
  FallThrough ft_s7_c1_r0(
    .io_a(ft_s7_c1_r0_io_a),
    .io_s(ft_s7_c1_r0_io_s)
  );
  wire ft_s8_c1_r0_io_a;
  wire ft_s8_c1_r0_io_s;
  FallThrough ft_s8_c1_r0(
    .io_a(ft_s8_c1_r0_io_a),
    .io_s(ft_s8_c1_r0_io_s)
  );
  wire ha_s0_c2_r0_io_a;
  wire ha_s0_c2_r0_io_b;
  wire ha_s0_c2_r0_io_s;
  wire ha_s0_c2_r0_io_co;
  HalfAdder ha_s0_c2_r0(
    .io_a(ha_s0_c2_r0_io_a),
    .io_b(ha_s0_c2_r0_io_b),
    .io_s(ha_s0_c2_r0_io_s),
    .io_co(ha_s0_c2_r0_io_co)
  );
  wire ft_s0_c2_r1_io_a;
  wire ft_s0_c2_r1_io_s;
  FallThrough ft_s0_c2_r1(
    .io_a(ft_s0_c2_r1_io_a),
    .io_s(ft_s0_c2_r1_io_s)
  );
  wire ha_s1_c2_r0_io_a;
  wire ha_s1_c2_r0_io_b;
  wire ha_s1_c2_r0_io_s;
  wire ha_s1_c2_r0_io_co;
  HalfAdder ha_s1_c2_r0(
    .io_a(ha_s1_c2_r0_io_a),
    .io_b(ha_s1_c2_r0_io_b),
    .io_s(ha_s1_c2_r0_io_s),
    .io_co(ha_s1_c2_r0_io_co)
  );
  wire ft_s1_c2_r1_io_a;
  wire ft_s1_c2_r1_io_s;
  FallThrough ft_s1_c2_r1(
    .io_a(ft_s1_c2_r1_io_a),
    .io_s(ft_s1_c2_r1_io_s)
  );
  wire ft_s2_c2_r0_io_a;
  wire ft_s2_c2_r0_io_s;
  FallThrough ft_s2_c2_r0(
    .io_a(ft_s2_c2_r0_io_a),
    .io_s(ft_s2_c2_r0_io_s)
  );
  wire ft_s2_c2_r1_io_a;
  wire ft_s2_c2_r1_io_s;
  FallThrough ft_s2_c2_r1(
    .io_a(ft_s2_c2_r1_io_a),
    .io_s(ft_s2_c2_r1_io_s)
  );
  wire ft_s3_c2_r0_io_a;
  wire ft_s3_c2_r0_io_s;
  FallThrough ft_s3_c2_r0(
    .io_a(ft_s3_c2_r0_io_a),
    .io_s(ft_s3_c2_r0_io_s)
  );
  wire ft_s3_c2_r1_io_a;
  wire ft_s3_c2_r1_io_s;
  FallThrough ft_s3_c2_r1(
    .io_a(ft_s3_c2_r1_io_a),
    .io_s(ft_s3_c2_r1_io_s)
  );
  wire ft_s4_c2_r0_io_a;
  wire ft_s4_c2_r0_io_s;
  FallThrough ft_s4_c2_r0(
    .io_a(ft_s4_c2_r0_io_a),
    .io_s(ft_s4_c2_r0_io_s)
  );
  wire ft_s4_c2_r1_io_a;
  wire ft_s4_c2_r1_io_s;
  FallThrough ft_s4_c2_r1(
    .io_a(ft_s4_c2_r1_io_a),
    .io_s(ft_s4_c2_r1_io_s)
  );
  wire ft_s5_c2_r0_io_a;
  wire ft_s5_c2_r0_io_s;
  FallThrough ft_s5_c2_r0(
    .io_a(ft_s5_c2_r0_io_a),
    .io_s(ft_s5_c2_r0_io_s)
  );
  wire ft_s5_c2_r1_io_a;
  wire ft_s5_c2_r1_io_s;
  FallThrough ft_s5_c2_r1(
    .io_a(ft_s5_c2_r1_io_a),
    .io_s(ft_s5_c2_r1_io_s)
  );
  wire ft_s6_c2_r0_io_a;
  wire ft_s6_c2_r0_io_s;
  FallThrough ft_s6_c2_r0(
    .io_a(ft_s6_c2_r0_io_a),
    .io_s(ft_s6_c2_r0_io_s)
  );
  wire ft_s6_c2_r1_io_a;
  wire ft_s6_c2_r1_io_s;
  FallThrough ft_s6_c2_r1(
    .io_a(ft_s6_c2_r1_io_a),
    .io_s(ft_s6_c2_r1_io_s)
  );
  wire ft_s7_c2_r0_io_a;
  wire ft_s7_c2_r0_io_s;
  FallThrough ft_s7_c2_r0(
    .io_a(ft_s7_c2_r0_io_a),
    .io_s(ft_s7_c2_r0_io_s)
  );
  wire ft_s7_c2_r1_io_a;
  wire ft_s7_c2_r1_io_s;
  FallThrough ft_s7_c2_r1(
    .io_a(ft_s7_c2_r1_io_a),
    .io_s(ft_s7_c2_r1_io_s)
  );
  wire ft_s8_c2_r0_io_a;
  wire ft_s8_c2_r0_io_s;
  FallThrough ft_s8_c2_r0(
    .io_a(ft_s8_c2_r0_io_a),
    .io_s(ft_s8_c2_r0_io_s)
  );
  wire ft_s8_c2_r1_io_a;
  wire ft_s8_c2_r1_io_s;
  FallThrough ft_s8_c2_r1(
    .io_a(ft_s8_c2_r1_io_a),
    .io_s(ft_s8_c2_r1_io_s)
  );
  wire fa_s0_c3_r0_io_a;
  wire fa_s0_c3_r0_io_b;
  wire fa_s0_c3_r0_io_ci;
  wire fa_s0_c3_r0_io_s;
  wire fa_s0_c3_r0_io_co;
  FullAdder fa_s0_c3_r0(
    .io_a(fa_s0_c3_r0_io_a),
    .io_b(fa_s0_c3_r0_io_b),
    .io_ci(fa_s0_c3_r0_io_ci),
    .io_s(fa_s0_c3_r0_io_s),
    .io_co(fa_s0_c3_r0_io_co)
  );
  wire ft_s0_c3_r1_io_a;
  wire ft_s0_c3_r1_io_s;
  FallThrough ft_s0_c3_r1(
    .io_a(ft_s0_c3_r1_io_a),
    .io_s(ft_s0_c3_r1_io_s)
  );
  wire fa_s1_c3_r0_io_a;
  wire fa_s1_c3_r0_io_b;
  wire fa_s1_c3_r0_io_ci;
  wire fa_s1_c3_r0_io_s;
  wire fa_s1_c3_r0_io_co;
  FullAdder fa_s1_c3_r0(
    .io_a(fa_s1_c3_r0_io_a),
    .io_b(fa_s1_c3_r0_io_b),
    .io_ci(fa_s1_c3_r0_io_ci),
    .io_s(fa_s1_c3_r0_io_s),
    .io_co(fa_s1_c3_r0_io_co)
  );
  wire ha_s2_c3_r0_io_a;
  wire ha_s2_c3_r0_io_b;
  wire ha_s2_c3_r0_io_s;
  wire ha_s2_c3_r0_io_co;
  HalfAdder ha_s2_c3_r0(
    .io_a(ha_s2_c3_r0_io_a),
    .io_b(ha_s2_c3_r0_io_b),
    .io_s(ha_s2_c3_r0_io_s),
    .io_co(ha_s2_c3_r0_io_co)
  );
  wire ft_s3_c3_r0_io_a;
  wire ft_s3_c3_r0_io_s;
  FallThrough ft_s3_c3_r0(
    .io_a(ft_s3_c3_r0_io_a),
    .io_s(ft_s3_c3_r0_io_s)
  );
  wire ft_s4_c3_r0_io_a;
  wire ft_s4_c3_r0_io_s;
  FallThrough ft_s4_c3_r0(
    .io_a(ft_s4_c3_r0_io_a),
    .io_s(ft_s4_c3_r0_io_s)
  );
  wire ft_s5_c3_r0_io_a;
  wire ft_s5_c3_r0_io_s;
  FallThrough ft_s5_c3_r0(
    .io_a(ft_s5_c3_r0_io_a),
    .io_s(ft_s5_c3_r0_io_s)
  );
  wire ft_s6_c3_r0_io_a;
  wire ft_s6_c3_r0_io_s;
  FallThrough ft_s6_c3_r0(
    .io_a(ft_s6_c3_r0_io_a),
    .io_s(ft_s6_c3_r0_io_s)
  );
  wire ft_s7_c3_r0_io_a;
  wire ft_s7_c3_r0_io_s;
  FallThrough ft_s7_c3_r0(
    .io_a(ft_s7_c3_r0_io_a),
    .io_s(ft_s7_c3_r0_io_s)
  );
  wire ft_s8_c3_r0_io_a;
  wire ft_s8_c3_r0_io_s;
  FallThrough ft_s8_c3_r0(
    .io_a(ft_s8_c3_r0_io_a),
    .io_s(ft_s8_c3_r0_io_s)
  );
  wire fa_s0_c4_r0_io_a;
  wire fa_s0_c4_r0_io_b;
  wire fa_s0_c4_r0_io_ci;
  wire fa_s0_c4_r0_io_s;
  wire fa_s0_c4_r0_io_co;
  FullAdder fa_s0_c4_r0(
    .io_a(fa_s0_c4_r0_io_a),
    .io_b(fa_s0_c4_r0_io_b),
    .io_ci(fa_s0_c4_r0_io_ci),
    .io_s(fa_s0_c4_r0_io_s),
    .io_co(fa_s0_c4_r0_io_co)
  );
  wire ft_s0_c4_r1_io_a;
  wire ft_s0_c4_r1_io_s;
  FallThrough ft_s0_c4_r1(
    .io_a(ft_s0_c4_r1_io_a),
    .io_s(ft_s0_c4_r1_io_s)
  );
  wire ft_s0_c4_r2_io_a;
  wire ft_s0_c4_r2_io_s;
  FallThrough ft_s0_c4_r2(
    .io_a(ft_s0_c4_r2_io_a),
    .io_s(ft_s0_c4_r2_io_s)
  );
  wire fa_s1_c4_r0_io_a;
  wire fa_s1_c4_r0_io_b;
  wire fa_s1_c4_r0_io_ci;
  wire fa_s1_c4_r0_io_s;
  wire fa_s1_c4_r0_io_co;
  FullAdder fa_s1_c4_r0(
    .io_a(fa_s1_c4_r0_io_a),
    .io_b(fa_s1_c4_r0_io_b),
    .io_ci(fa_s1_c4_r0_io_ci),
    .io_s(fa_s1_c4_r0_io_s),
    .io_co(fa_s1_c4_r0_io_co)
  );
  wire ft_s1_c4_r1_io_a;
  wire ft_s1_c4_r1_io_s;
  FallThrough ft_s1_c4_r1(
    .io_a(ft_s1_c4_r1_io_a),
    .io_s(ft_s1_c4_r1_io_s)
  );
  wire fa_s2_c4_r0_io_a;
  wire fa_s2_c4_r0_io_b;
  wire fa_s2_c4_r0_io_ci;
  wire fa_s2_c4_r0_io_s;
  wire fa_s2_c4_r0_io_co;
  FullAdder fa_s2_c4_r0(
    .io_a(fa_s2_c4_r0_io_a),
    .io_b(fa_s2_c4_r0_io_b),
    .io_ci(fa_s2_c4_r0_io_ci),
    .io_s(fa_s2_c4_r0_io_s),
    .io_co(fa_s2_c4_r0_io_co)
  );
  wire ft_s3_c4_r0_io_a;
  wire ft_s3_c4_r0_io_s;
  FallThrough ft_s3_c4_r0(
    .io_a(ft_s3_c4_r0_io_a),
    .io_s(ft_s3_c4_r0_io_s)
  );
  wire ft_s3_c4_r1_io_a;
  wire ft_s3_c4_r1_io_s;
  FallThrough ft_s3_c4_r1(
    .io_a(ft_s3_c4_r1_io_a),
    .io_s(ft_s3_c4_r1_io_s)
  );
  wire ft_s4_c4_r0_io_a;
  wire ft_s4_c4_r0_io_s;
  FallThrough ft_s4_c4_r0(
    .io_a(ft_s4_c4_r0_io_a),
    .io_s(ft_s4_c4_r0_io_s)
  );
  wire ft_s4_c4_r1_io_a;
  wire ft_s4_c4_r1_io_s;
  FallThrough ft_s4_c4_r1(
    .io_a(ft_s4_c4_r1_io_a),
    .io_s(ft_s4_c4_r1_io_s)
  );
  wire ft_s5_c4_r0_io_a;
  wire ft_s5_c4_r0_io_s;
  FallThrough ft_s5_c4_r0(
    .io_a(ft_s5_c4_r0_io_a),
    .io_s(ft_s5_c4_r0_io_s)
  );
  wire ft_s5_c4_r1_io_a;
  wire ft_s5_c4_r1_io_s;
  FallThrough ft_s5_c4_r1(
    .io_a(ft_s5_c4_r1_io_a),
    .io_s(ft_s5_c4_r1_io_s)
  );
  wire ft_s6_c4_r0_io_a;
  wire ft_s6_c4_r0_io_s;
  FallThrough ft_s6_c4_r0(
    .io_a(ft_s6_c4_r0_io_a),
    .io_s(ft_s6_c4_r0_io_s)
  );
  wire ft_s6_c4_r1_io_a;
  wire ft_s6_c4_r1_io_s;
  FallThrough ft_s6_c4_r1(
    .io_a(ft_s6_c4_r1_io_a),
    .io_s(ft_s6_c4_r1_io_s)
  );
  wire ft_s7_c4_r0_io_a;
  wire ft_s7_c4_r0_io_s;
  FallThrough ft_s7_c4_r0(
    .io_a(ft_s7_c4_r0_io_a),
    .io_s(ft_s7_c4_r0_io_s)
  );
  wire ft_s7_c4_r1_io_a;
  wire ft_s7_c4_r1_io_s;
  FallThrough ft_s7_c4_r1(
    .io_a(ft_s7_c4_r1_io_a),
    .io_s(ft_s7_c4_r1_io_s)
  );
  wire ft_s8_c4_r0_io_a;
  wire ft_s8_c4_r0_io_s;
  FallThrough ft_s8_c4_r0(
    .io_a(ft_s8_c4_r0_io_a),
    .io_s(ft_s8_c4_r0_io_s)
  );
  wire ft_s8_c4_r1_io_a;
  wire ft_s8_c4_r1_io_s;
  FallThrough ft_s8_c4_r1(
    .io_a(ft_s8_c4_r1_io_a),
    .io_s(ft_s8_c4_r1_io_s)
  );
  wire fa_s0_c5_r0_io_a;
  wire fa_s0_c5_r0_io_b;
  wire fa_s0_c5_r0_io_ci;
  wire fa_s0_c5_r0_io_s;
  wire fa_s0_c5_r0_io_co;
  FullAdder fa_s0_c5_r0(
    .io_a(fa_s0_c5_r0_io_a),
    .io_b(fa_s0_c5_r0_io_b),
    .io_ci(fa_s0_c5_r0_io_ci),
    .io_s(fa_s0_c5_r0_io_s),
    .io_co(fa_s0_c5_r0_io_co)
  );
  wire fa_s0_c5_r1_io_a;
  wire fa_s0_c5_r1_io_b;
  wire fa_s0_c5_r1_io_ci;
  wire fa_s0_c5_r1_io_s;
  wire fa_s0_c5_r1_io_co;
  FullAdder fa_s0_c5_r1(
    .io_a(fa_s0_c5_r1_io_a),
    .io_b(fa_s0_c5_r1_io_b),
    .io_ci(fa_s0_c5_r1_io_ci),
    .io_s(fa_s0_c5_r1_io_s),
    .io_co(fa_s0_c5_r1_io_co)
  );
  wire fa_s1_c5_r0_io_a;
  wire fa_s1_c5_r0_io_b;
  wire fa_s1_c5_r0_io_ci;
  wire fa_s1_c5_r0_io_s;
  wire fa_s1_c5_r0_io_co;
  FullAdder fa_s1_c5_r0(
    .io_a(fa_s1_c5_r0_io_a),
    .io_b(fa_s1_c5_r0_io_b),
    .io_ci(fa_s1_c5_r0_io_ci),
    .io_s(fa_s1_c5_r0_io_s),
    .io_co(fa_s1_c5_r0_io_co)
  );
  wire ft_s2_c5_r0_io_a;
  wire ft_s2_c5_r0_io_s;
  FallThrough ft_s2_c5_r0(
    .io_a(ft_s2_c5_r0_io_a),
    .io_s(ft_s2_c5_r0_io_s)
  );
  wire ft_s2_c5_r1_io_a;
  wire ft_s2_c5_r1_io_s;
  FallThrough ft_s2_c5_r1(
    .io_a(ft_s2_c5_r1_io_a),
    .io_s(ft_s2_c5_r1_io_s)
  );
  wire fa_s3_c5_r0_io_a;
  wire fa_s3_c5_r0_io_b;
  wire fa_s3_c5_r0_io_ci;
  wire fa_s3_c5_r0_io_s;
  wire fa_s3_c5_r0_io_co;
  FullAdder fa_s3_c5_r0(
    .io_a(fa_s3_c5_r0_io_a),
    .io_b(fa_s3_c5_r0_io_b),
    .io_ci(fa_s3_c5_r0_io_ci),
    .io_s(fa_s3_c5_r0_io_s),
    .io_co(fa_s3_c5_r0_io_co)
  );
  wire ft_s4_c5_r0_io_a;
  wire ft_s4_c5_r0_io_s;
  FallThrough ft_s4_c5_r0(
    .io_a(ft_s4_c5_r0_io_a),
    .io_s(ft_s4_c5_r0_io_s)
  );
  wire ft_s5_c5_r0_io_a;
  wire ft_s5_c5_r0_io_s;
  FallThrough ft_s5_c5_r0(
    .io_a(ft_s5_c5_r0_io_a),
    .io_s(ft_s5_c5_r0_io_s)
  );
  wire ft_s6_c5_r0_io_a;
  wire ft_s6_c5_r0_io_s;
  FallThrough ft_s6_c5_r0(
    .io_a(ft_s6_c5_r0_io_a),
    .io_s(ft_s6_c5_r0_io_s)
  );
  wire ft_s7_c5_r0_io_a;
  wire ft_s7_c5_r0_io_s;
  FallThrough ft_s7_c5_r0(
    .io_a(ft_s7_c5_r0_io_a),
    .io_s(ft_s7_c5_r0_io_s)
  );
  wire ft_s8_c5_r0_io_a;
  wire ft_s8_c5_r0_io_s;
  FallThrough ft_s8_c5_r0(
    .io_a(ft_s8_c5_r0_io_a),
    .io_s(ft_s8_c5_r0_io_s)
  );
  wire fa_s0_c6_r0_io_a;
  wire fa_s0_c6_r0_io_b;
  wire fa_s0_c6_r0_io_ci;
  wire fa_s0_c6_r0_io_s;
  wire fa_s0_c6_r0_io_co;
  FullAdder fa_s0_c6_r0(
    .io_a(fa_s0_c6_r0_io_a),
    .io_b(fa_s0_c6_r0_io_b),
    .io_ci(fa_s0_c6_r0_io_ci),
    .io_s(fa_s0_c6_r0_io_s),
    .io_co(fa_s0_c6_r0_io_co)
  );
  wire fa_s0_c6_r1_io_a;
  wire fa_s0_c6_r1_io_b;
  wire fa_s0_c6_r1_io_ci;
  wire fa_s0_c6_r1_io_s;
  wire fa_s0_c6_r1_io_co;
  FullAdder fa_s0_c6_r1(
    .io_a(fa_s0_c6_r1_io_a),
    .io_b(fa_s0_c6_r1_io_b),
    .io_ci(fa_s0_c6_r1_io_ci),
    .io_s(fa_s0_c6_r1_io_s),
    .io_co(fa_s0_c6_r1_io_co)
  );
  wire ft_s0_c6_r2_io_a;
  wire ft_s0_c6_r2_io_s;
  FallThrough ft_s0_c6_r2(
    .io_a(ft_s0_c6_r2_io_a),
    .io_s(ft_s0_c6_r2_io_s)
  );
  wire fa_s1_c6_r0_io_a;
  wire fa_s1_c6_r0_io_b;
  wire fa_s1_c6_r0_io_ci;
  wire fa_s1_c6_r0_io_s;
  wire fa_s1_c6_r0_io_co;
  FullAdder fa_s1_c6_r0(
    .io_a(fa_s1_c6_r0_io_a),
    .io_b(fa_s1_c6_r0_io_b),
    .io_ci(fa_s1_c6_r0_io_ci),
    .io_s(fa_s1_c6_r0_io_s),
    .io_co(fa_s1_c6_r0_io_co)
  );
  wire ha_s1_c6_r1_io_a;
  wire ha_s1_c6_r1_io_b;
  wire ha_s1_c6_r1_io_s;
  wire ha_s1_c6_r1_io_co;
  HalfAdder ha_s1_c6_r1(
    .io_a(ha_s1_c6_r1_io_a),
    .io_b(ha_s1_c6_r1_io_b),
    .io_s(ha_s1_c6_r1_io_s),
    .io_co(ha_s1_c6_r1_io_co)
  );
  wire fa_s2_c6_r0_io_a;
  wire fa_s2_c6_r0_io_b;
  wire fa_s2_c6_r0_io_ci;
  wire fa_s2_c6_r0_io_s;
  wire fa_s2_c6_r0_io_co;
  FullAdder fa_s2_c6_r0(
    .io_a(fa_s2_c6_r0_io_a),
    .io_b(fa_s2_c6_r0_io_b),
    .io_ci(fa_s2_c6_r0_io_ci),
    .io_s(fa_s2_c6_r0_io_s),
    .io_co(fa_s2_c6_r0_io_co)
  );
  wire ft_s3_c6_r0_io_a;
  wire ft_s3_c6_r0_io_s;
  FallThrough ft_s3_c6_r0(
    .io_a(ft_s3_c6_r0_io_a),
    .io_s(ft_s3_c6_r0_io_s)
  );
  wire ft_s4_c6_r0_io_a;
  wire ft_s4_c6_r0_io_s;
  FallThrough ft_s4_c6_r0(
    .io_a(ft_s4_c6_r0_io_a),
    .io_s(ft_s4_c6_r0_io_s)
  );
  wire ft_s4_c6_r1_io_a;
  wire ft_s4_c6_r1_io_s;
  FallThrough ft_s4_c6_r1(
    .io_a(ft_s4_c6_r1_io_a),
    .io_s(ft_s4_c6_r1_io_s)
  );
  wire ft_s5_c6_r0_io_a;
  wire ft_s5_c6_r0_io_s;
  FallThrough ft_s5_c6_r0(
    .io_a(ft_s5_c6_r0_io_a),
    .io_s(ft_s5_c6_r0_io_s)
  );
  wire ft_s5_c6_r1_io_a;
  wire ft_s5_c6_r1_io_s;
  FallThrough ft_s5_c6_r1(
    .io_a(ft_s5_c6_r1_io_a),
    .io_s(ft_s5_c6_r1_io_s)
  );
  wire ft_s6_c6_r0_io_a;
  wire ft_s6_c6_r0_io_s;
  FallThrough ft_s6_c6_r0(
    .io_a(ft_s6_c6_r0_io_a),
    .io_s(ft_s6_c6_r0_io_s)
  );
  wire ft_s6_c6_r1_io_a;
  wire ft_s6_c6_r1_io_s;
  FallThrough ft_s6_c6_r1(
    .io_a(ft_s6_c6_r1_io_a),
    .io_s(ft_s6_c6_r1_io_s)
  );
  wire ft_s7_c6_r0_io_a;
  wire ft_s7_c6_r0_io_s;
  FallThrough ft_s7_c6_r0(
    .io_a(ft_s7_c6_r0_io_a),
    .io_s(ft_s7_c6_r0_io_s)
  );
  wire ft_s7_c6_r1_io_a;
  wire ft_s7_c6_r1_io_s;
  FallThrough ft_s7_c6_r1(
    .io_a(ft_s7_c6_r1_io_a),
    .io_s(ft_s7_c6_r1_io_s)
  );
  wire ft_s8_c6_r0_io_a;
  wire ft_s8_c6_r0_io_s;
  FallThrough ft_s8_c6_r0(
    .io_a(ft_s8_c6_r0_io_a),
    .io_s(ft_s8_c6_r0_io_s)
  );
  wire ft_s8_c6_r1_io_a;
  wire ft_s8_c6_r1_io_s;
  FallThrough ft_s8_c6_r1(
    .io_a(ft_s8_c6_r1_io_a),
    .io_s(ft_s8_c6_r1_io_s)
  );
  wire fa_s0_c7_r0_io_a;
  wire fa_s0_c7_r0_io_b;
  wire fa_s0_c7_r0_io_ci;
  wire fa_s0_c7_r0_io_s;
  wire fa_s0_c7_r0_io_co;
  FullAdder fa_s0_c7_r0(
    .io_a(fa_s0_c7_r0_io_a),
    .io_b(fa_s0_c7_r0_io_b),
    .io_ci(fa_s0_c7_r0_io_ci),
    .io_s(fa_s0_c7_r0_io_s),
    .io_co(fa_s0_c7_r0_io_co)
  );
  wire fa_s0_c7_r1_io_a;
  wire fa_s0_c7_r1_io_b;
  wire fa_s0_c7_r1_io_ci;
  wire fa_s0_c7_r1_io_s;
  wire fa_s0_c7_r1_io_co;
  FullAdder fa_s0_c7_r1(
    .io_a(fa_s0_c7_r1_io_a),
    .io_b(fa_s0_c7_r1_io_b),
    .io_ci(fa_s0_c7_r1_io_ci),
    .io_s(fa_s0_c7_r1_io_s),
    .io_co(fa_s0_c7_r1_io_co)
  );
  wire ft_s0_c7_r2_io_a;
  wire ft_s0_c7_r2_io_s;
  FallThrough ft_s0_c7_r2(
    .io_a(ft_s0_c7_r2_io_a),
    .io_s(ft_s0_c7_r2_io_s)
  );
  wire ft_s0_c7_r3_io_a;
  wire ft_s0_c7_r3_io_s;
  FallThrough ft_s0_c7_r3(
    .io_a(ft_s0_c7_r3_io_a),
    .io_s(ft_s0_c7_r3_io_s)
  );
  wire fa_s1_c7_r0_io_a;
  wire fa_s1_c7_r0_io_b;
  wire fa_s1_c7_r0_io_ci;
  wire fa_s1_c7_r0_io_s;
  wire fa_s1_c7_r0_io_co;
  FullAdder fa_s1_c7_r0(
    .io_a(fa_s1_c7_r0_io_a),
    .io_b(fa_s1_c7_r0_io_b),
    .io_ci(fa_s1_c7_r0_io_ci),
    .io_s(fa_s1_c7_r0_io_s),
    .io_co(fa_s1_c7_r0_io_co)
  );
  wire fa_s1_c7_r1_io_a;
  wire fa_s1_c7_r1_io_b;
  wire fa_s1_c7_r1_io_ci;
  wire fa_s1_c7_r1_io_s;
  wire fa_s1_c7_r1_io_co;
  FullAdder fa_s1_c7_r1(
    .io_a(fa_s1_c7_r1_io_a),
    .io_b(fa_s1_c7_r1_io_b),
    .io_ci(fa_s1_c7_r1_io_ci),
    .io_s(fa_s1_c7_r1_io_s),
    .io_co(fa_s1_c7_r1_io_co)
  );
  wire fa_s2_c7_r0_io_a;
  wire fa_s2_c7_r0_io_b;
  wire fa_s2_c7_r0_io_ci;
  wire fa_s2_c7_r0_io_s;
  wire fa_s2_c7_r0_io_co;
  FullAdder fa_s2_c7_r0(
    .io_a(fa_s2_c7_r0_io_a),
    .io_b(fa_s2_c7_r0_io_b),
    .io_ci(fa_s2_c7_r0_io_ci),
    .io_s(fa_s2_c7_r0_io_s),
    .io_co(fa_s2_c7_r0_io_co)
  );
  wire ft_s2_c7_r1_io_a;
  wire ft_s2_c7_r1_io_s;
  FallThrough ft_s2_c7_r1(
    .io_a(ft_s2_c7_r1_io_a),
    .io_s(ft_s2_c7_r1_io_s)
  );
  wire fa_s3_c7_r0_io_a;
  wire fa_s3_c7_r0_io_b;
  wire fa_s3_c7_r0_io_ci;
  wire fa_s3_c7_r0_io_s;
  wire fa_s3_c7_r0_io_co;
  FullAdder fa_s3_c7_r0(
    .io_a(fa_s3_c7_r0_io_a),
    .io_b(fa_s3_c7_r0_io_b),
    .io_ci(fa_s3_c7_r0_io_ci),
    .io_s(fa_s3_c7_r0_io_s),
    .io_co(fa_s3_c7_r0_io_co)
  );
  wire ft_s4_c7_r0_io_a;
  wire ft_s4_c7_r0_io_s;
  FallThrough ft_s4_c7_r0(
    .io_a(ft_s4_c7_r0_io_a),
    .io_s(ft_s4_c7_r0_io_s)
  );
  wire ft_s5_c7_r0_io_a;
  wire ft_s5_c7_r0_io_s;
  FallThrough ft_s5_c7_r0(
    .io_a(ft_s5_c7_r0_io_a),
    .io_s(ft_s5_c7_r0_io_s)
  );
  wire ft_s6_c7_r0_io_a;
  wire ft_s6_c7_r0_io_s;
  FallThrough ft_s6_c7_r0(
    .io_a(ft_s6_c7_r0_io_a),
    .io_s(ft_s6_c7_r0_io_s)
  );
  wire ft_s7_c7_r0_io_a;
  wire ft_s7_c7_r0_io_s;
  FallThrough ft_s7_c7_r0(
    .io_a(ft_s7_c7_r0_io_a),
    .io_s(ft_s7_c7_r0_io_s)
  );
  wire ft_s8_c7_r0_io_a;
  wire ft_s8_c7_r0_io_s;
  FallThrough ft_s8_c7_r0(
    .io_a(ft_s8_c7_r0_io_a),
    .io_s(ft_s8_c7_r0_io_s)
  );
  wire fa_s0_c8_r0_io_a;
  wire fa_s0_c8_r0_io_b;
  wire fa_s0_c8_r0_io_ci;
  wire fa_s0_c8_r0_io_s;
  wire fa_s0_c8_r0_io_co;
  FullAdder fa_s0_c8_r0(
    .io_a(fa_s0_c8_r0_io_a),
    .io_b(fa_s0_c8_r0_io_b),
    .io_ci(fa_s0_c8_r0_io_ci),
    .io_s(fa_s0_c8_r0_io_s),
    .io_co(fa_s0_c8_r0_io_co)
  );
  wire fa_s0_c8_r1_io_a;
  wire fa_s0_c8_r1_io_b;
  wire fa_s0_c8_r1_io_ci;
  wire fa_s0_c8_r1_io_s;
  wire fa_s0_c8_r1_io_co;
  FullAdder fa_s0_c8_r1(
    .io_a(fa_s0_c8_r1_io_a),
    .io_b(fa_s0_c8_r1_io_b),
    .io_ci(fa_s0_c8_r1_io_ci),
    .io_s(fa_s0_c8_r1_io_s),
    .io_co(fa_s0_c8_r1_io_co)
  );
  wire fa_s0_c8_r2_io_a;
  wire fa_s0_c8_r2_io_b;
  wire fa_s0_c8_r2_io_ci;
  wire fa_s0_c8_r2_io_s;
  wire fa_s0_c8_r2_io_co;
  FullAdder fa_s0_c8_r2(
    .io_a(fa_s0_c8_r2_io_a),
    .io_b(fa_s0_c8_r2_io_b),
    .io_ci(fa_s0_c8_r2_io_ci),
    .io_s(fa_s0_c8_r2_io_s),
    .io_co(fa_s0_c8_r2_io_co)
  );
  wire fa_s1_c8_r0_io_a;
  wire fa_s1_c8_r0_io_b;
  wire fa_s1_c8_r0_io_ci;
  wire fa_s1_c8_r0_io_s;
  wire fa_s1_c8_r0_io_co;
  FullAdder fa_s1_c8_r0(
    .io_a(fa_s1_c8_r0_io_a),
    .io_b(fa_s1_c8_r0_io_b),
    .io_ci(fa_s1_c8_r0_io_ci),
    .io_s(fa_s1_c8_r0_io_s),
    .io_co(fa_s1_c8_r0_io_co)
  );
  wire ha_s1_c8_r1_io_a;
  wire ha_s1_c8_r1_io_b;
  wire ha_s1_c8_r1_io_s;
  wire ha_s1_c8_r1_io_co;
  HalfAdder ha_s1_c8_r1(
    .io_a(ha_s1_c8_r1_io_a),
    .io_b(ha_s1_c8_r1_io_b),
    .io_s(ha_s1_c8_r1_io_s),
    .io_co(ha_s1_c8_r1_io_co)
  );
  wire fa_s2_c8_r0_io_a;
  wire fa_s2_c8_r0_io_b;
  wire fa_s2_c8_r0_io_ci;
  wire fa_s2_c8_r0_io_s;
  wire fa_s2_c8_r0_io_co;
  FullAdder fa_s2_c8_r0(
    .io_a(fa_s2_c8_r0_io_a),
    .io_b(fa_s2_c8_r0_io_b),
    .io_ci(fa_s2_c8_r0_io_ci),
    .io_s(fa_s2_c8_r0_io_s),
    .io_co(fa_s2_c8_r0_io_co)
  );
  wire ft_s2_c8_r1_io_a;
  wire ft_s2_c8_r1_io_s;
  FallThrough ft_s2_c8_r1(
    .io_a(ft_s2_c8_r1_io_a),
    .io_s(ft_s2_c8_r1_io_s)
  );
  wire fa_s3_c8_r0_io_a;
  wire fa_s3_c8_r0_io_b;
  wire fa_s3_c8_r0_io_ci;
  wire fa_s3_c8_r0_io_s;
  wire fa_s3_c8_r0_io_co;
  FullAdder fa_s3_c8_r0(
    .io_a(fa_s3_c8_r0_io_a),
    .io_b(fa_s3_c8_r0_io_b),
    .io_ci(fa_s3_c8_r0_io_ci),
    .io_s(fa_s3_c8_r0_io_s),
    .io_co(fa_s3_c8_r0_io_co)
  );
  wire ft_s4_c8_r0_io_a;
  wire ft_s4_c8_r0_io_s;
  FallThrough ft_s4_c8_r0(
    .io_a(ft_s4_c8_r0_io_a),
    .io_s(ft_s4_c8_r0_io_s)
  );
  wire ft_s4_c8_r1_io_a;
  wire ft_s4_c8_r1_io_s;
  FallThrough ft_s4_c8_r1(
    .io_a(ft_s4_c8_r1_io_a),
    .io_s(ft_s4_c8_r1_io_s)
  );
  wire ft_s5_c8_r0_io_a;
  wire ft_s5_c8_r0_io_s;
  FallThrough ft_s5_c8_r0(
    .io_a(ft_s5_c8_r0_io_a),
    .io_s(ft_s5_c8_r0_io_s)
  );
  wire ft_s5_c8_r1_io_a;
  wire ft_s5_c8_r1_io_s;
  FallThrough ft_s5_c8_r1(
    .io_a(ft_s5_c8_r1_io_a),
    .io_s(ft_s5_c8_r1_io_s)
  );
  wire ft_s6_c8_r0_io_a;
  wire ft_s6_c8_r0_io_s;
  FallThrough ft_s6_c8_r0(
    .io_a(ft_s6_c8_r0_io_a),
    .io_s(ft_s6_c8_r0_io_s)
  );
  wire ft_s6_c8_r1_io_a;
  wire ft_s6_c8_r1_io_s;
  FallThrough ft_s6_c8_r1(
    .io_a(ft_s6_c8_r1_io_a),
    .io_s(ft_s6_c8_r1_io_s)
  );
  wire ft_s7_c8_r0_io_a;
  wire ft_s7_c8_r0_io_s;
  FallThrough ft_s7_c8_r0(
    .io_a(ft_s7_c8_r0_io_a),
    .io_s(ft_s7_c8_r0_io_s)
  );
  wire ft_s7_c8_r1_io_a;
  wire ft_s7_c8_r1_io_s;
  FallThrough ft_s7_c8_r1(
    .io_a(ft_s7_c8_r1_io_a),
    .io_s(ft_s7_c8_r1_io_s)
  );
  wire ft_s8_c8_r0_io_a;
  wire ft_s8_c8_r0_io_s;
  FallThrough ft_s8_c8_r0(
    .io_a(ft_s8_c8_r0_io_a),
    .io_s(ft_s8_c8_r0_io_s)
  );
  wire ft_s8_c8_r1_io_a;
  wire ft_s8_c8_r1_io_s;
  FallThrough ft_s8_c8_r1(
    .io_a(ft_s8_c8_r1_io_a),
    .io_s(ft_s8_c8_r1_io_s)
  );
  wire fa_s0_c9_r0_io_a;
  wire fa_s0_c9_r0_io_b;
  wire fa_s0_c9_r0_io_ci;
  wire fa_s0_c9_r0_io_s;
  wire fa_s0_c9_r0_io_co;
  FullAdder fa_s0_c9_r0(
    .io_a(fa_s0_c9_r0_io_a),
    .io_b(fa_s0_c9_r0_io_b),
    .io_ci(fa_s0_c9_r0_io_ci),
    .io_s(fa_s0_c9_r0_io_s),
    .io_co(fa_s0_c9_r0_io_co)
  );
  wire fa_s0_c9_r1_io_a;
  wire fa_s0_c9_r1_io_b;
  wire fa_s0_c9_r1_io_ci;
  wire fa_s0_c9_r1_io_s;
  wire fa_s0_c9_r1_io_co;
  FullAdder fa_s0_c9_r1(
    .io_a(fa_s0_c9_r1_io_a),
    .io_b(fa_s0_c9_r1_io_b),
    .io_ci(fa_s0_c9_r1_io_ci),
    .io_s(fa_s0_c9_r1_io_s),
    .io_co(fa_s0_c9_r1_io_co)
  );
  wire fa_s0_c9_r2_io_a;
  wire fa_s0_c9_r2_io_b;
  wire fa_s0_c9_r2_io_ci;
  wire fa_s0_c9_r2_io_s;
  wire fa_s0_c9_r2_io_co;
  FullAdder fa_s0_c9_r2(
    .io_a(fa_s0_c9_r2_io_a),
    .io_b(fa_s0_c9_r2_io_b),
    .io_ci(fa_s0_c9_r2_io_ci),
    .io_s(fa_s0_c9_r2_io_s),
    .io_co(fa_s0_c9_r2_io_co)
  );
  wire ft_s0_c9_r3_io_a;
  wire ft_s0_c9_r3_io_s;
  FallThrough ft_s0_c9_r3(
    .io_a(ft_s0_c9_r3_io_a),
    .io_s(ft_s0_c9_r3_io_s)
  );
  wire fa_s1_c9_r0_io_a;
  wire fa_s1_c9_r0_io_b;
  wire fa_s1_c9_r0_io_ci;
  wire fa_s1_c9_r0_io_s;
  wire fa_s1_c9_r0_io_co;
  FullAdder fa_s1_c9_r0(
    .io_a(fa_s1_c9_r0_io_a),
    .io_b(fa_s1_c9_r0_io_b),
    .io_ci(fa_s1_c9_r0_io_ci),
    .io_s(fa_s1_c9_r0_io_s),
    .io_co(fa_s1_c9_r0_io_co)
  );
  wire fa_s1_c9_r1_io_a;
  wire fa_s1_c9_r1_io_b;
  wire fa_s1_c9_r1_io_ci;
  wire fa_s1_c9_r1_io_s;
  wire fa_s1_c9_r1_io_co;
  FullAdder fa_s1_c9_r1(
    .io_a(fa_s1_c9_r1_io_a),
    .io_b(fa_s1_c9_r1_io_b),
    .io_ci(fa_s1_c9_r1_io_ci),
    .io_s(fa_s1_c9_r1_io_s),
    .io_co(fa_s1_c9_r1_io_co)
  );
  wire ft_s1_c9_r2_io_a;
  wire ft_s1_c9_r2_io_s;
  FallThrough ft_s1_c9_r2(
    .io_a(ft_s1_c9_r2_io_a),
    .io_s(ft_s1_c9_r2_io_s)
  );
  wire ha_s2_c9_r0_io_a;
  wire ha_s2_c9_r0_io_b;
  wire ha_s2_c9_r0_io_s;
  wire ha_s2_c9_r0_io_co;
  HalfAdder ha_s2_c9_r0(
    .io_a(ha_s2_c9_r0_io_a),
    .io_b(ha_s2_c9_r0_io_b),
    .io_s(ha_s2_c9_r0_io_s),
    .io_co(ha_s2_c9_r0_io_co)
  );
  wire ha_s2_c9_r1_io_a;
  wire ha_s2_c9_r1_io_b;
  wire ha_s2_c9_r1_io_s;
  wire ha_s2_c9_r1_io_co;
  HalfAdder ha_s2_c9_r1(
    .io_a(ha_s2_c9_r1_io_a),
    .io_b(ha_s2_c9_r1_io_b),
    .io_s(ha_s2_c9_r1_io_s),
    .io_co(ha_s2_c9_r1_io_co)
  );
  wire ft_s2_c9_r2_io_a;
  wire ft_s2_c9_r2_io_s;
  FallThrough ft_s2_c9_r2(
    .io_a(ft_s2_c9_r2_io_a),
    .io_s(ft_s2_c9_r2_io_s)
  );
  wire ha_s3_c9_r0_io_a;
  wire ha_s3_c9_r0_io_b;
  wire ha_s3_c9_r0_io_s;
  wire ha_s3_c9_r0_io_co;
  HalfAdder ha_s3_c9_r0(
    .io_a(ha_s3_c9_r0_io_a),
    .io_b(ha_s3_c9_r0_io_b),
    .io_s(ha_s3_c9_r0_io_s),
    .io_co(ha_s3_c9_r0_io_co)
  );
  wire ft_s3_c9_r1_io_a;
  wire ft_s3_c9_r1_io_s;
  FallThrough ft_s3_c9_r1(
    .io_a(ft_s3_c9_r1_io_a),
    .io_s(ft_s3_c9_r1_io_s)
  );
  wire ft_s3_c9_r2_io_a;
  wire ft_s3_c9_r2_io_s;
  FallThrough ft_s3_c9_r2(
    .io_a(ft_s3_c9_r2_io_a),
    .io_s(ft_s3_c9_r2_io_s)
  );
  wire ha_s4_c9_r0_io_a;
  wire ha_s4_c9_r0_io_b;
  wire ha_s4_c9_r0_io_s;
  wire ha_s4_c9_r0_io_co;
  HalfAdder ha_s4_c9_r0(
    .io_a(ha_s4_c9_r0_io_a),
    .io_b(ha_s4_c9_r0_io_b),
    .io_s(ha_s4_c9_r0_io_s),
    .io_co(ha_s4_c9_r0_io_co)
  );
  wire ft_s4_c9_r1_io_a;
  wire ft_s4_c9_r1_io_s;
  FallThrough ft_s4_c9_r1(
    .io_a(ft_s4_c9_r1_io_a),
    .io_s(ft_s4_c9_r1_io_s)
  );
  wire ft_s4_c9_r2_io_a;
  wire ft_s4_c9_r2_io_s;
  FallThrough ft_s4_c9_r2(
    .io_a(ft_s4_c9_r2_io_a),
    .io_s(ft_s4_c9_r2_io_s)
  );
  wire fa_s5_c9_r0_io_a;
  wire fa_s5_c9_r0_io_b;
  wire fa_s5_c9_r0_io_ci;
  wire fa_s5_c9_r0_io_s;
  wire fa_s5_c9_r0_io_co;
  FullAdder fa_s5_c9_r0(
    .io_a(fa_s5_c9_r0_io_a),
    .io_b(fa_s5_c9_r0_io_b),
    .io_ci(fa_s5_c9_r0_io_ci),
    .io_s(fa_s5_c9_r0_io_s),
    .io_co(fa_s5_c9_r0_io_co)
  );
  wire ft_s6_c9_r0_io_a;
  wire ft_s6_c9_r0_io_s;
  FallThrough ft_s6_c9_r0(
    .io_a(ft_s6_c9_r0_io_a),
    .io_s(ft_s6_c9_r0_io_s)
  );
  wire ft_s7_c9_r0_io_a;
  wire ft_s7_c9_r0_io_s;
  FallThrough ft_s7_c9_r0(
    .io_a(ft_s7_c9_r0_io_a),
    .io_s(ft_s7_c9_r0_io_s)
  );
  wire ft_s8_c9_r0_io_a;
  wire ft_s8_c9_r0_io_s;
  FallThrough ft_s8_c9_r0(
    .io_a(ft_s8_c9_r0_io_a),
    .io_s(ft_s8_c9_r0_io_s)
  );
  wire fa_s0_c10_r0_io_a;
  wire fa_s0_c10_r0_io_b;
  wire fa_s0_c10_r0_io_ci;
  wire fa_s0_c10_r0_io_s;
  wire fa_s0_c10_r0_io_co;
  FullAdder fa_s0_c10_r0(
    .io_a(fa_s0_c10_r0_io_a),
    .io_b(fa_s0_c10_r0_io_b),
    .io_ci(fa_s0_c10_r0_io_ci),
    .io_s(fa_s0_c10_r0_io_s),
    .io_co(fa_s0_c10_r0_io_co)
  );
  wire fa_s0_c10_r1_io_a;
  wire fa_s0_c10_r1_io_b;
  wire fa_s0_c10_r1_io_ci;
  wire fa_s0_c10_r1_io_s;
  wire fa_s0_c10_r1_io_co;
  FullAdder fa_s0_c10_r1(
    .io_a(fa_s0_c10_r1_io_a),
    .io_b(fa_s0_c10_r1_io_b),
    .io_ci(fa_s0_c10_r1_io_ci),
    .io_s(fa_s0_c10_r1_io_s),
    .io_co(fa_s0_c10_r1_io_co)
  );
  wire fa_s0_c10_r2_io_a;
  wire fa_s0_c10_r2_io_b;
  wire fa_s0_c10_r2_io_ci;
  wire fa_s0_c10_r2_io_s;
  wire fa_s0_c10_r2_io_co;
  FullAdder fa_s0_c10_r2(
    .io_a(fa_s0_c10_r2_io_a),
    .io_b(fa_s0_c10_r2_io_b),
    .io_ci(fa_s0_c10_r2_io_ci),
    .io_s(fa_s0_c10_r2_io_s),
    .io_co(fa_s0_c10_r2_io_co)
  );
  wire ft_s0_c10_r3_io_a;
  wire ft_s0_c10_r3_io_s;
  FallThrough ft_s0_c10_r3(
    .io_a(ft_s0_c10_r3_io_a),
    .io_s(ft_s0_c10_r3_io_s)
  );
  wire ft_s0_c10_r4_io_a;
  wire ft_s0_c10_r4_io_s;
  FallThrough ft_s0_c10_r4(
    .io_a(ft_s0_c10_r4_io_a),
    .io_s(ft_s0_c10_r4_io_s)
  );
  wire fa_s1_c10_r0_io_a;
  wire fa_s1_c10_r0_io_b;
  wire fa_s1_c10_r0_io_ci;
  wire fa_s1_c10_r0_io_s;
  wire fa_s1_c10_r0_io_co;
  FullAdder fa_s1_c10_r0(
    .io_a(fa_s1_c10_r0_io_a),
    .io_b(fa_s1_c10_r0_io_b),
    .io_ci(fa_s1_c10_r0_io_ci),
    .io_s(fa_s1_c10_r0_io_s),
    .io_co(fa_s1_c10_r0_io_co)
  );
  wire fa_s1_c10_r1_io_a;
  wire fa_s1_c10_r1_io_b;
  wire fa_s1_c10_r1_io_ci;
  wire fa_s1_c10_r1_io_s;
  wire fa_s1_c10_r1_io_co;
  FullAdder fa_s1_c10_r1(
    .io_a(fa_s1_c10_r1_io_a),
    .io_b(fa_s1_c10_r1_io_b),
    .io_ci(fa_s1_c10_r1_io_ci),
    .io_s(fa_s1_c10_r1_io_s),
    .io_co(fa_s1_c10_r1_io_co)
  );
  wire ft_s1_c10_r2_io_a;
  wire ft_s1_c10_r2_io_s;
  FallThrough ft_s1_c10_r2(
    .io_a(ft_s1_c10_r2_io_a),
    .io_s(ft_s1_c10_r2_io_s)
  );
  wire ft_s1_c10_r3_io_a;
  wire ft_s1_c10_r3_io_s;
  FallThrough ft_s1_c10_r3(
    .io_a(ft_s1_c10_r3_io_a),
    .io_s(ft_s1_c10_r3_io_s)
  );
  wire fa_s2_c10_r0_io_a;
  wire fa_s2_c10_r0_io_b;
  wire fa_s2_c10_r0_io_ci;
  wire fa_s2_c10_r0_io_s;
  wire fa_s2_c10_r0_io_co;
  FullAdder fa_s2_c10_r0(
    .io_a(fa_s2_c10_r0_io_a),
    .io_b(fa_s2_c10_r0_io_b),
    .io_ci(fa_s2_c10_r0_io_ci),
    .io_s(fa_s2_c10_r0_io_s),
    .io_co(fa_s2_c10_r0_io_co)
  );
  wire fa_s2_c10_r1_io_a;
  wire fa_s2_c10_r1_io_b;
  wire fa_s2_c10_r1_io_ci;
  wire fa_s2_c10_r1_io_s;
  wire fa_s2_c10_r1_io_co;
  FullAdder fa_s2_c10_r1(
    .io_a(fa_s2_c10_r1_io_a),
    .io_b(fa_s2_c10_r1_io_b),
    .io_ci(fa_s2_c10_r1_io_ci),
    .io_s(fa_s2_c10_r1_io_s),
    .io_co(fa_s2_c10_r1_io_co)
  );
  wire fa_s3_c10_r0_io_a;
  wire fa_s3_c10_r0_io_b;
  wire fa_s3_c10_r0_io_ci;
  wire fa_s3_c10_r0_io_s;
  wire fa_s3_c10_r0_io_co;
  FullAdder fa_s3_c10_r0(
    .io_a(fa_s3_c10_r0_io_a),
    .io_b(fa_s3_c10_r0_io_b),
    .io_ci(fa_s3_c10_r0_io_ci),
    .io_s(fa_s3_c10_r0_io_s),
    .io_co(fa_s3_c10_r0_io_co)
  );
  wire ft_s3_c10_r1_io_a;
  wire ft_s3_c10_r1_io_s;
  FallThrough ft_s3_c10_r1(
    .io_a(ft_s3_c10_r1_io_a),
    .io_s(ft_s3_c10_r1_io_s)
  );
  wire fa_s4_c10_r0_io_a;
  wire fa_s4_c10_r0_io_b;
  wire fa_s4_c10_r0_io_ci;
  wire fa_s4_c10_r0_io_s;
  wire fa_s4_c10_r0_io_co;
  FullAdder fa_s4_c10_r0(
    .io_a(fa_s4_c10_r0_io_a),
    .io_b(fa_s4_c10_r0_io_b),
    .io_ci(fa_s4_c10_r0_io_ci),
    .io_s(fa_s4_c10_r0_io_s),
    .io_co(fa_s4_c10_r0_io_co)
  );
  wire ft_s5_c10_r0_io_a;
  wire ft_s5_c10_r0_io_s;
  FallThrough ft_s5_c10_r0(
    .io_a(ft_s5_c10_r0_io_a),
    .io_s(ft_s5_c10_r0_io_s)
  );
  wire ft_s5_c10_r1_io_a;
  wire ft_s5_c10_r1_io_s;
  FallThrough ft_s5_c10_r1(
    .io_a(ft_s5_c10_r1_io_a),
    .io_s(ft_s5_c10_r1_io_s)
  );
  wire fa_s6_c10_r0_io_a;
  wire fa_s6_c10_r0_io_b;
  wire fa_s6_c10_r0_io_ci;
  wire fa_s6_c10_r0_io_s;
  wire fa_s6_c10_r0_io_co;
  FullAdder fa_s6_c10_r0(
    .io_a(fa_s6_c10_r0_io_a),
    .io_b(fa_s6_c10_r0_io_b),
    .io_ci(fa_s6_c10_r0_io_ci),
    .io_s(fa_s6_c10_r0_io_s),
    .io_co(fa_s6_c10_r0_io_co)
  );
  wire ft_s7_c10_r0_io_a;
  wire ft_s7_c10_r0_io_s;
  FallThrough ft_s7_c10_r0(
    .io_a(ft_s7_c10_r0_io_a),
    .io_s(ft_s7_c10_r0_io_s)
  );
  wire ft_s8_c10_r0_io_a;
  wire ft_s8_c10_r0_io_s;
  FallThrough ft_s8_c10_r0(
    .io_a(ft_s8_c10_r0_io_a),
    .io_s(ft_s8_c10_r0_io_s)
  );
  wire fa_s0_c11_r0_io_a;
  wire fa_s0_c11_r0_io_b;
  wire fa_s0_c11_r0_io_ci;
  wire fa_s0_c11_r0_io_s;
  wire fa_s0_c11_r0_io_co;
  FullAdder fa_s0_c11_r0(
    .io_a(fa_s0_c11_r0_io_a),
    .io_b(fa_s0_c11_r0_io_b),
    .io_ci(fa_s0_c11_r0_io_ci),
    .io_s(fa_s0_c11_r0_io_s),
    .io_co(fa_s0_c11_r0_io_co)
  );
  wire fa_s0_c11_r1_io_a;
  wire fa_s0_c11_r1_io_b;
  wire fa_s0_c11_r1_io_ci;
  wire fa_s0_c11_r1_io_s;
  wire fa_s0_c11_r1_io_co;
  FullAdder fa_s0_c11_r1(
    .io_a(fa_s0_c11_r1_io_a),
    .io_b(fa_s0_c11_r1_io_b),
    .io_ci(fa_s0_c11_r1_io_ci),
    .io_s(fa_s0_c11_r1_io_s),
    .io_co(fa_s0_c11_r1_io_co)
  );
  wire fa_s0_c11_r2_io_a;
  wire fa_s0_c11_r2_io_b;
  wire fa_s0_c11_r2_io_ci;
  wire fa_s0_c11_r2_io_s;
  wire fa_s0_c11_r2_io_co;
  FullAdder fa_s0_c11_r2(
    .io_a(fa_s0_c11_r2_io_a),
    .io_b(fa_s0_c11_r2_io_b),
    .io_ci(fa_s0_c11_r2_io_ci),
    .io_s(fa_s0_c11_r2_io_s),
    .io_co(fa_s0_c11_r2_io_co)
  );
  wire fa_s0_c11_r3_io_a;
  wire fa_s0_c11_r3_io_b;
  wire fa_s0_c11_r3_io_ci;
  wire fa_s0_c11_r3_io_s;
  wire fa_s0_c11_r3_io_co;
  FullAdder fa_s0_c11_r3(
    .io_a(fa_s0_c11_r3_io_a),
    .io_b(fa_s0_c11_r3_io_b),
    .io_ci(fa_s0_c11_r3_io_ci),
    .io_s(fa_s0_c11_r3_io_s),
    .io_co(fa_s0_c11_r3_io_co)
  );
  wire fa_s1_c11_r0_io_a;
  wire fa_s1_c11_r0_io_b;
  wire fa_s1_c11_r0_io_ci;
  wire fa_s1_c11_r0_io_s;
  wire fa_s1_c11_r0_io_co;
  FullAdder fa_s1_c11_r0(
    .io_a(fa_s1_c11_r0_io_a),
    .io_b(fa_s1_c11_r0_io_b),
    .io_ci(fa_s1_c11_r0_io_ci),
    .io_s(fa_s1_c11_r0_io_s),
    .io_co(fa_s1_c11_r0_io_co)
  );
  wire fa_s1_c11_r1_io_a;
  wire fa_s1_c11_r1_io_b;
  wire fa_s1_c11_r1_io_ci;
  wire fa_s1_c11_r1_io_s;
  wire fa_s1_c11_r1_io_co;
  FullAdder fa_s1_c11_r1(
    .io_a(fa_s1_c11_r1_io_a),
    .io_b(fa_s1_c11_r1_io_b),
    .io_ci(fa_s1_c11_r1_io_ci),
    .io_s(fa_s1_c11_r1_io_s),
    .io_co(fa_s1_c11_r1_io_co)
  );
  wire ft_s1_c11_r2_io_a;
  wire ft_s1_c11_r2_io_s;
  FallThrough ft_s1_c11_r2(
    .io_a(ft_s1_c11_r2_io_a),
    .io_s(ft_s1_c11_r2_io_s)
  );
  wire fa_s2_c11_r0_io_a;
  wire fa_s2_c11_r0_io_b;
  wire fa_s2_c11_r0_io_ci;
  wire fa_s2_c11_r0_io_s;
  wire fa_s2_c11_r0_io_co;
  FullAdder fa_s2_c11_r0(
    .io_a(fa_s2_c11_r0_io_a),
    .io_b(fa_s2_c11_r0_io_b),
    .io_ci(fa_s2_c11_r0_io_ci),
    .io_s(fa_s2_c11_r0_io_s),
    .io_co(fa_s2_c11_r0_io_co)
  );
  wire ha_s2_c11_r1_io_a;
  wire ha_s2_c11_r1_io_b;
  wire ha_s2_c11_r1_io_s;
  wire ha_s2_c11_r1_io_co;
  HalfAdder ha_s2_c11_r1(
    .io_a(ha_s2_c11_r1_io_a),
    .io_b(ha_s2_c11_r1_io_b),
    .io_s(ha_s2_c11_r1_io_s),
    .io_co(ha_s2_c11_r1_io_co)
  );
  wire fa_s3_c11_r0_io_a;
  wire fa_s3_c11_r0_io_b;
  wire fa_s3_c11_r0_io_ci;
  wire fa_s3_c11_r0_io_s;
  wire fa_s3_c11_r0_io_co;
  FullAdder fa_s3_c11_r0(
    .io_a(fa_s3_c11_r0_io_a),
    .io_b(fa_s3_c11_r0_io_b),
    .io_ci(fa_s3_c11_r0_io_ci),
    .io_s(fa_s3_c11_r0_io_s),
    .io_co(fa_s3_c11_r0_io_co)
  );
  wire ft_s3_c11_r1_io_a;
  wire ft_s3_c11_r1_io_s;
  FallThrough ft_s3_c11_r1(
    .io_a(ft_s3_c11_r1_io_a),
    .io_s(ft_s3_c11_r1_io_s)
  );
  wire ha_s4_c11_r0_io_a;
  wire ha_s4_c11_r0_io_b;
  wire ha_s4_c11_r0_io_s;
  wire ha_s4_c11_r0_io_co;
  HalfAdder ha_s4_c11_r0(
    .io_a(ha_s4_c11_r0_io_a),
    .io_b(ha_s4_c11_r0_io_b),
    .io_s(ha_s4_c11_r0_io_s),
    .io_co(ha_s4_c11_r0_io_co)
  );
  wire ft_s4_c11_r1_io_a;
  wire ft_s4_c11_r1_io_s;
  FallThrough ft_s4_c11_r1(
    .io_a(ft_s4_c11_r1_io_a),
    .io_s(ft_s4_c11_r1_io_s)
  );
  wire ha_s5_c11_r0_io_a;
  wire ha_s5_c11_r0_io_b;
  wire ha_s5_c11_r0_io_s;
  wire ha_s5_c11_r0_io_co;
  HalfAdder ha_s5_c11_r0(
    .io_a(ha_s5_c11_r0_io_a),
    .io_b(ha_s5_c11_r0_io_b),
    .io_s(ha_s5_c11_r0_io_s),
    .io_co(ha_s5_c11_r0_io_co)
  );
  wire ft_s5_c11_r1_io_a;
  wire ft_s5_c11_r1_io_s;
  FallThrough ft_s5_c11_r1(
    .io_a(ft_s5_c11_r1_io_a),
    .io_s(ft_s5_c11_r1_io_s)
  );
  wire ha_s6_c11_r0_io_a;
  wire ha_s6_c11_r0_io_b;
  wire ha_s6_c11_r0_io_s;
  wire ha_s6_c11_r0_io_co;
  HalfAdder ha_s6_c11_r0(
    .io_a(ha_s6_c11_r0_io_a),
    .io_b(ha_s6_c11_r0_io_b),
    .io_s(ha_s6_c11_r0_io_s),
    .io_co(ha_s6_c11_r0_io_co)
  );
  wire ft_s7_c11_r0_io_a;
  wire ft_s7_c11_r0_io_s;
  FallThrough ft_s7_c11_r0(
    .io_a(ft_s7_c11_r0_io_a),
    .io_s(ft_s7_c11_r0_io_s)
  );
  wire ft_s7_c11_r1_io_a;
  wire ft_s7_c11_r1_io_s;
  FallThrough ft_s7_c11_r1(
    .io_a(ft_s7_c11_r1_io_a),
    .io_s(ft_s7_c11_r1_io_s)
  );
  wire ft_s8_c11_r0_io_a;
  wire ft_s8_c11_r0_io_s;
  FallThrough ft_s8_c11_r0(
    .io_a(ft_s8_c11_r0_io_a),
    .io_s(ft_s8_c11_r0_io_s)
  );
  wire ft_s8_c11_r1_io_a;
  wire ft_s8_c11_r1_io_s;
  FallThrough ft_s8_c11_r1(
    .io_a(ft_s8_c11_r1_io_a),
    .io_s(ft_s8_c11_r1_io_s)
  );
  wire fa_s0_c12_r0_io_a;
  wire fa_s0_c12_r0_io_b;
  wire fa_s0_c12_r0_io_ci;
  wire fa_s0_c12_r0_io_s;
  wire fa_s0_c12_r0_io_co;
  FullAdder fa_s0_c12_r0(
    .io_a(fa_s0_c12_r0_io_a),
    .io_b(fa_s0_c12_r0_io_b),
    .io_ci(fa_s0_c12_r0_io_ci),
    .io_s(fa_s0_c12_r0_io_s),
    .io_co(fa_s0_c12_r0_io_co)
  );
  wire fa_s0_c12_r1_io_a;
  wire fa_s0_c12_r1_io_b;
  wire fa_s0_c12_r1_io_ci;
  wire fa_s0_c12_r1_io_s;
  wire fa_s0_c12_r1_io_co;
  FullAdder fa_s0_c12_r1(
    .io_a(fa_s0_c12_r1_io_a),
    .io_b(fa_s0_c12_r1_io_b),
    .io_ci(fa_s0_c12_r1_io_ci),
    .io_s(fa_s0_c12_r1_io_s),
    .io_co(fa_s0_c12_r1_io_co)
  );
  wire fa_s0_c12_r2_io_a;
  wire fa_s0_c12_r2_io_b;
  wire fa_s0_c12_r2_io_ci;
  wire fa_s0_c12_r2_io_s;
  wire fa_s0_c12_r2_io_co;
  FullAdder fa_s0_c12_r2(
    .io_a(fa_s0_c12_r2_io_a),
    .io_b(fa_s0_c12_r2_io_b),
    .io_ci(fa_s0_c12_r2_io_ci),
    .io_s(fa_s0_c12_r2_io_s),
    .io_co(fa_s0_c12_r2_io_co)
  );
  wire fa_s0_c12_r3_io_a;
  wire fa_s0_c12_r3_io_b;
  wire fa_s0_c12_r3_io_ci;
  wire fa_s0_c12_r3_io_s;
  wire fa_s0_c12_r3_io_co;
  FullAdder fa_s0_c12_r3(
    .io_a(fa_s0_c12_r3_io_a),
    .io_b(fa_s0_c12_r3_io_b),
    .io_ci(fa_s0_c12_r3_io_ci),
    .io_s(fa_s0_c12_r3_io_s),
    .io_co(fa_s0_c12_r3_io_co)
  );
  wire ft_s0_c12_r4_io_a;
  wire ft_s0_c12_r4_io_s;
  FallThrough ft_s0_c12_r4(
    .io_a(ft_s0_c12_r4_io_a),
    .io_s(ft_s0_c12_r4_io_s)
  );
  wire fa_s1_c12_r0_io_a;
  wire fa_s1_c12_r0_io_b;
  wire fa_s1_c12_r0_io_ci;
  wire fa_s1_c12_r0_io_s;
  wire fa_s1_c12_r0_io_co;
  FullAdder fa_s1_c12_r0(
    .io_a(fa_s1_c12_r0_io_a),
    .io_b(fa_s1_c12_r0_io_b),
    .io_ci(fa_s1_c12_r0_io_ci),
    .io_s(fa_s1_c12_r0_io_s),
    .io_co(fa_s1_c12_r0_io_co)
  );
  wire fa_s1_c12_r1_io_a;
  wire fa_s1_c12_r1_io_b;
  wire fa_s1_c12_r1_io_ci;
  wire fa_s1_c12_r1_io_s;
  wire fa_s1_c12_r1_io_co;
  FullAdder fa_s1_c12_r1(
    .io_a(fa_s1_c12_r1_io_a),
    .io_b(fa_s1_c12_r1_io_b),
    .io_ci(fa_s1_c12_r1_io_ci),
    .io_s(fa_s1_c12_r1_io_s),
    .io_co(fa_s1_c12_r1_io_co)
  );
  wire fa_s1_c12_r2_io_a;
  wire fa_s1_c12_r2_io_b;
  wire fa_s1_c12_r2_io_ci;
  wire fa_s1_c12_r2_io_s;
  wire fa_s1_c12_r2_io_co;
  FullAdder fa_s1_c12_r2(
    .io_a(fa_s1_c12_r2_io_a),
    .io_b(fa_s1_c12_r2_io_b),
    .io_ci(fa_s1_c12_r2_io_ci),
    .io_s(fa_s1_c12_r2_io_s),
    .io_co(fa_s1_c12_r2_io_co)
  );
  wire fa_s2_c12_r0_io_a;
  wire fa_s2_c12_r0_io_b;
  wire fa_s2_c12_r0_io_ci;
  wire fa_s2_c12_r0_io_s;
  wire fa_s2_c12_r0_io_co;
  FullAdder fa_s2_c12_r0(
    .io_a(fa_s2_c12_r0_io_a),
    .io_b(fa_s2_c12_r0_io_b),
    .io_ci(fa_s2_c12_r0_io_ci),
    .io_s(fa_s2_c12_r0_io_s),
    .io_co(fa_s2_c12_r0_io_co)
  );
  wire ft_s2_c12_r1_io_a;
  wire ft_s2_c12_r1_io_s;
  FallThrough ft_s2_c12_r1(
    .io_a(ft_s2_c12_r1_io_a),
    .io_s(ft_s2_c12_r1_io_s)
  );
  wire ft_s2_c12_r2_io_a;
  wire ft_s2_c12_r2_io_s;
  FallThrough ft_s2_c12_r2(
    .io_a(ft_s2_c12_r2_io_a),
    .io_s(ft_s2_c12_r2_io_s)
  );
  wire fa_s3_c12_r0_io_a;
  wire fa_s3_c12_r0_io_b;
  wire fa_s3_c12_r0_io_ci;
  wire fa_s3_c12_r0_io_s;
  wire fa_s3_c12_r0_io_co;
  FullAdder fa_s3_c12_r0(
    .io_a(fa_s3_c12_r0_io_a),
    .io_b(fa_s3_c12_r0_io_b),
    .io_ci(fa_s3_c12_r0_io_ci),
    .io_s(fa_s3_c12_r0_io_s),
    .io_co(fa_s3_c12_r0_io_co)
  );
  wire ft_s3_c12_r1_io_a;
  wire ft_s3_c12_r1_io_s;
  FallThrough ft_s3_c12_r1(
    .io_a(ft_s3_c12_r1_io_a),
    .io_s(ft_s3_c12_r1_io_s)
  );
  wire ft_s3_c12_r2_io_a;
  wire ft_s3_c12_r2_io_s;
  FallThrough ft_s3_c12_r2(
    .io_a(ft_s3_c12_r2_io_a),
    .io_s(ft_s3_c12_r2_io_s)
  );
  wire fa_s4_c12_r0_io_a;
  wire fa_s4_c12_r0_io_b;
  wire fa_s4_c12_r0_io_ci;
  wire fa_s4_c12_r0_io_s;
  wire fa_s4_c12_r0_io_co;
  FullAdder fa_s4_c12_r0(
    .io_a(fa_s4_c12_r0_io_a),
    .io_b(fa_s4_c12_r0_io_b),
    .io_ci(fa_s4_c12_r0_io_ci),
    .io_s(fa_s4_c12_r0_io_s),
    .io_co(fa_s4_c12_r0_io_co)
  );
  wire ft_s4_c12_r1_io_a;
  wire ft_s4_c12_r1_io_s;
  FallThrough ft_s4_c12_r1(
    .io_a(ft_s4_c12_r1_io_a),
    .io_s(ft_s4_c12_r1_io_s)
  );
  wire fa_s5_c12_r0_io_a;
  wire fa_s5_c12_r0_io_b;
  wire fa_s5_c12_r0_io_ci;
  wire fa_s5_c12_r0_io_s;
  wire fa_s5_c12_r0_io_co;
  FullAdder fa_s5_c12_r0(
    .io_a(fa_s5_c12_r0_io_a),
    .io_b(fa_s5_c12_r0_io_b),
    .io_ci(fa_s5_c12_r0_io_ci),
    .io_s(fa_s5_c12_r0_io_s),
    .io_co(fa_s5_c12_r0_io_co)
  );
  wire ft_s6_c12_r0_io_a;
  wire ft_s6_c12_r0_io_s;
  FallThrough ft_s6_c12_r0(
    .io_a(ft_s6_c12_r0_io_a),
    .io_s(ft_s6_c12_r0_io_s)
  );
  wire ft_s6_c12_r1_io_a;
  wire ft_s6_c12_r1_io_s;
  FallThrough ft_s6_c12_r1(
    .io_a(ft_s6_c12_r1_io_a),
    .io_s(ft_s6_c12_r1_io_s)
  );
  wire fa_s7_c12_r0_io_a;
  wire fa_s7_c12_r0_io_b;
  wire fa_s7_c12_r0_io_ci;
  wire fa_s7_c12_r0_io_s;
  wire fa_s7_c12_r0_io_co;
  FullAdder fa_s7_c12_r0(
    .io_a(fa_s7_c12_r0_io_a),
    .io_b(fa_s7_c12_r0_io_b),
    .io_ci(fa_s7_c12_r0_io_ci),
    .io_s(fa_s7_c12_r0_io_s),
    .io_co(fa_s7_c12_r0_io_co)
  );
  wire ft_s8_c12_r0_io_a;
  wire ft_s8_c12_r0_io_s;
  FallThrough ft_s8_c12_r0(
    .io_a(ft_s8_c12_r0_io_a),
    .io_s(ft_s8_c12_r0_io_s)
  );
  wire fa_s0_c13_r0_io_a;
  wire fa_s0_c13_r0_io_b;
  wire fa_s0_c13_r0_io_ci;
  wire fa_s0_c13_r0_io_s;
  wire fa_s0_c13_r0_io_co;
  FullAdder fa_s0_c13_r0(
    .io_a(fa_s0_c13_r0_io_a),
    .io_b(fa_s0_c13_r0_io_b),
    .io_ci(fa_s0_c13_r0_io_ci),
    .io_s(fa_s0_c13_r0_io_s),
    .io_co(fa_s0_c13_r0_io_co)
  );
  wire fa_s0_c13_r1_io_a;
  wire fa_s0_c13_r1_io_b;
  wire fa_s0_c13_r1_io_ci;
  wire fa_s0_c13_r1_io_s;
  wire fa_s0_c13_r1_io_co;
  FullAdder fa_s0_c13_r1(
    .io_a(fa_s0_c13_r1_io_a),
    .io_b(fa_s0_c13_r1_io_b),
    .io_ci(fa_s0_c13_r1_io_ci),
    .io_s(fa_s0_c13_r1_io_s),
    .io_co(fa_s0_c13_r1_io_co)
  );
  wire fa_s0_c13_r2_io_a;
  wire fa_s0_c13_r2_io_b;
  wire fa_s0_c13_r2_io_ci;
  wire fa_s0_c13_r2_io_s;
  wire fa_s0_c13_r2_io_co;
  FullAdder fa_s0_c13_r2(
    .io_a(fa_s0_c13_r2_io_a),
    .io_b(fa_s0_c13_r2_io_b),
    .io_ci(fa_s0_c13_r2_io_ci),
    .io_s(fa_s0_c13_r2_io_s),
    .io_co(fa_s0_c13_r2_io_co)
  );
  wire fa_s0_c13_r3_io_a;
  wire fa_s0_c13_r3_io_b;
  wire fa_s0_c13_r3_io_ci;
  wire fa_s0_c13_r3_io_s;
  wire fa_s0_c13_r3_io_co;
  FullAdder fa_s0_c13_r3(
    .io_a(fa_s0_c13_r3_io_a),
    .io_b(fa_s0_c13_r3_io_b),
    .io_ci(fa_s0_c13_r3_io_ci),
    .io_s(fa_s0_c13_r3_io_s),
    .io_co(fa_s0_c13_r3_io_co)
  );
  wire ft_s0_c13_r4_io_a;
  wire ft_s0_c13_r4_io_s;
  FallThrough ft_s0_c13_r4(
    .io_a(ft_s0_c13_r4_io_a),
    .io_s(ft_s0_c13_r4_io_s)
  );
  wire ft_s0_c13_r5_io_a;
  wire ft_s0_c13_r5_io_s;
  FallThrough ft_s0_c13_r5(
    .io_a(ft_s0_c13_r5_io_a),
    .io_s(ft_s0_c13_r5_io_s)
  );
  wire fa_s1_c13_r0_io_a;
  wire fa_s1_c13_r0_io_b;
  wire fa_s1_c13_r0_io_ci;
  wire fa_s1_c13_r0_io_s;
  wire fa_s1_c13_r0_io_co;
  FullAdder fa_s1_c13_r0(
    .io_a(fa_s1_c13_r0_io_a),
    .io_b(fa_s1_c13_r0_io_b),
    .io_ci(fa_s1_c13_r0_io_ci),
    .io_s(fa_s1_c13_r0_io_s),
    .io_co(fa_s1_c13_r0_io_co)
  );
  wire fa_s1_c13_r1_io_a;
  wire fa_s1_c13_r1_io_b;
  wire fa_s1_c13_r1_io_ci;
  wire fa_s1_c13_r1_io_s;
  wire fa_s1_c13_r1_io_co;
  FullAdder fa_s1_c13_r1(
    .io_a(fa_s1_c13_r1_io_a),
    .io_b(fa_s1_c13_r1_io_b),
    .io_ci(fa_s1_c13_r1_io_ci),
    .io_s(fa_s1_c13_r1_io_s),
    .io_co(fa_s1_c13_r1_io_co)
  );
  wire fa_s1_c13_r2_io_a;
  wire fa_s1_c13_r2_io_b;
  wire fa_s1_c13_r2_io_ci;
  wire fa_s1_c13_r2_io_s;
  wire fa_s1_c13_r2_io_co;
  FullAdder fa_s1_c13_r2(
    .io_a(fa_s1_c13_r2_io_a),
    .io_b(fa_s1_c13_r2_io_b),
    .io_ci(fa_s1_c13_r2_io_ci),
    .io_s(fa_s1_c13_r2_io_s),
    .io_co(fa_s1_c13_r2_io_co)
  );
  wire ft_s1_c13_r3_io_a;
  wire ft_s1_c13_r3_io_s;
  FallThrough ft_s1_c13_r3(
    .io_a(ft_s1_c13_r3_io_a),
    .io_s(ft_s1_c13_r3_io_s)
  );
  wire fa_s2_c13_r0_io_a;
  wire fa_s2_c13_r0_io_b;
  wire fa_s2_c13_r0_io_ci;
  wire fa_s2_c13_r0_io_s;
  wire fa_s2_c13_r0_io_co;
  FullAdder fa_s2_c13_r0(
    .io_a(fa_s2_c13_r0_io_a),
    .io_b(fa_s2_c13_r0_io_b),
    .io_ci(fa_s2_c13_r0_io_ci),
    .io_s(fa_s2_c13_r0_io_s),
    .io_co(fa_s2_c13_r0_io_co)
  );
  wire fa_s2_c13_r1_io_a;
  wire fa_s2_c13_r1_io_b;
  wire fa_s2_c13_r1_io_ci;
  wire fa_s2_c13_r1_io_s;
  wire fa_s2_c13_r1_io_co;
  FullAdder fa_s2_c13_r1(
    .io_a(fa_s2_c13_r1_io_a),
    .io_b(fa_s2_c13_r1_io_b),
    .io_ci(fa_s2_c13_r1_io_ci),
    .io_s(fa_s2_c13_r1_io_s),
    .io_co(fa_s2_c13_r1_io_co)
  );
  wire ft_s2_c13_r2_io_a;
  wire ft_s2_c13_r2_io_s;
  FallThrough ft_s2_c13_r2(
    .io_a(ft_s2_c13_r2_io_a),
    .io_s(ft_s2_c13_r2_io_s)
  );
  wire fa_s3_c13_r0_io_a;
  wire fa_s3_c13_r0_io_b;
  wire fa_s3_c13_r0_io_ci;
  wire fa_s3_c13_r0_io_s;
  wire fa_s3_c13_r0_io_co;
  FullAdder fa_s3_c13_r0(
    .io_a(fa_s3_c13_r0_io_a),
    .io_b(fa_s3_c13_r0_io_b),
    .io_ci(fa_s3_c13_r0_io_ci),
    .io_s(fa_s3_c13_r0_io_s),
    .io_co(fa_s3_c13_r0_io_co)
  );
  wire ft_s3_c13_r1_io_a;
  wire ft_s3_c13_r1_io_s;
  FallThrough ft_s3_c13_r1(
    .io_a(ft_s3_c13_r1_io_a),
    .io_s(ft_s3_c13_r1_io_s)
  );
  wire fa_s4_c13_r0_io_a;
  wire fa_s4_c13_r0_io_b;
  wire fa_s4_c13_r0_io_ci;
  wire fa_s4_c13_r0_io_s;
  wire fa_s4_c13_r0_io_co;
  FullAdder fa_s4_c13_r0(
    .io_a(fa_s4_c13_r0_io_a),
    .io_b(fa_s4_c13_r0_io_b),
    .io_ci(fa_s4_c13_r0_io_ci),
    .io_s(fa_s4_c13_r0_io_s),
    .io_co(fa_s4_c13_r0_io_co)
  );
  wire ft_s5_c13_r0_io_a;
  wire ft_s5_c13_r0_io_s;
  FallThrough ft_s5_c13_r0(
    .io_a(ft_s5_c13_r0_io_a),
    .io_s(ft_s5_c13_r0_io_s)
  );
  wire ft_s5_c13_r1_io_a;
  wire ft_s5_c13_r1_io_s;
  FallThrough ft_s5_c13_r1(
    .io_a(ft_s5_c13_r1_io_a),
    .io_s(ft_s5_c13_r1_io_s)
  );
  wire fa_s6_c13_r0_io_a;
  wire fa_s6_c13_r0_io_b;
  wire fa_s6_c13_r0_io_ci;
  wire fa_s6_c13_r0_io_s;
  wire fa_s6_c13_r0_io_co;
  FullAdder fa_s6_c13_r0(
    .io_a(fa_s6_c13_r0_io_a),
    .io_b(fa_s6_c13_r0_io_b),
    .io_ci(fa_s6_c13_r0_io_ci),
    .io_s(fa_s6_c13_r0_io_s),
    .io_co(fa_s6_c13_r0_io_co)
  );
  wire ft_s7_c13_r0_io_a;
  wire ft_s7_c13_r0_io_s;
  FallThrough ft_s7_c13_r0(
    .io_a(ft_s7_c13_r0_io_a),
    .io_s(ft_s7_c13_r0_io_s)
  );
  wire ft_s8_c13_r0_io_a;
  wire ft_s8_c13_r0_io_s;
  FallThrough ft_s8_c13_r0(
    .io_a(ft_s8_c13_r0_io_a),
    .io_s(ft_s8_c13_r0_io_s)
  );
  wire ft_s8_c13_r1_io_a;
  wire ft_s8_c13_r1_io_s;
  FallThrough ft_s8_c13_r1(
    .io_a(ft_s8_c13_r1_io_a),
    .io_s(ft_s8_c13_r1_io_s)
  );
  wire fa_s0_c14_r0_io_a;
  wire fa_s0_c14_r0_io_b;
  wire fa_s0_c14_r0_io_ci;
  wire fa_s0_c14_r0_io_s;
  wire fa_s0_c14_r0_io_co;
  FullAdder fa_s0_c14_r0(
    .io_a(fa_s0_c14_r0_io_a),
    .io_b(fa_s0_c14_r0_io_b),
    .io_ci(fa_s0_c14_r0_io_ci),
    .io_s(fa_s0_c14_r0_io_s),
    .io_co(fa_s0_c14_r0_io_co)
  );
  wire fa_s0_c14_r1_io_a;
  wire fa_s0_c14_r1_io_b;
  wire fa_s0_c14_r1_io_ci;
  wire fa_s0_c14_r1_io_s;
  wire fa_s0_c14_r1_io_co;
  FullAdder fa_s0_c14_r1(
    .io_a(fa_s0_c14_r1_io_a),
    .io_b(fa_s0_c14_r1_io_b),
    .io_ci(fa_s0_c14_r1_io_ci),
    .io_s(fa_s0_c14_r1_io_s),
    .io_co(fa_s0_c14_r1_io_co)
  );
  wire fa_s0_c14_r2_io_a;
  wire fa_s0_c14_r2_io_b;
  wire fa_s0_c14_r2_io_ci;
  wire fa_s0_c14_r2_io_s;
  wire fa_s0_c14_r2_io_co;
  FullAdder fa_s0_c14_r2(
    .io_a(fa_s0_c14_r2_io_a),
    .io_b(fa_s0_c14_r2_io_b),
    .io_ci(fa_s0_c14_r2_io_ci),
    .io_s(fa_s0_c14_r2_io_s),
    .io_co(fa_s0_c14_r2_io_co)
  );
  wire fa_s0_c14_r3_io_a;
  wire fa_s0_c14_r3_io_b;
  wire fa_s0_c14_r3_io_ci;
  wire fa_s0_c14_r3_io_s;
  wire fa_s0_c14_r3_io_co;
  FullAdder fa_s0_c14_r3(
    .io_a(fa_s0_c14_r3_io_a),
    .io_b(fa_s0_c14_r3_io_b),
    .io_ci(fa_s0_c14_r3_io_ci),
    .io_s(fa_s0_c14_r3_io_s),
    .io_co(fa_s0_c14_r3_io_co)
  );
  wire fa_s0_c14_r4_io_a;
  wire fa_s0_c14_r4_io_b;
  wire fa_s0_c14_r4_io_ci;
  wire fa_s0_c14_r4_io_s;
  wire fa_s0_c14_r4_io_co;
  FullAdder fa_s0_c14_r4(
    .io_a(fa_s0_c14_r4_io_a),
    .io_b(fa_s0_c14_r4_io_b),
    .io_ci(fa_s0_c14_r4_io_ci),
    .io_s(fa_s0_c14_r4_io_s),
    .io_co(fa_s0_c14_r4_io_co)
  );
  wire fa_s1_c14_r0_io_a;
  wire fa_s1_c14_r0_io_b;
  wire fa_s1_c14_r0_io_ci;
  wire fa_s1_c14_r0_io_s;
  wire fa_s1_c14_r0_io_co;
  FullAdder fa_s1_c14_r0(
    .io_a(fa_s1_c14_r0_io_a),
    .io_b(fa_s1_c14_r0_io_b),
    .io_ci(fa_s1_c14_r0_io_ci),
    .io_s(fa_s1_c14_r0_io_s),
    .io_co(fa_s1_c14_r0_io_co)
  );
  wire fa_s1_c14_r1_io_a;
  wire fa_s1_c14_r1_io_b;
  wire fa_s1_c14_r1_io_ci;
  wire fa_s1_c14_r1_io_s;
  wire fa_s1_c14_r1_io_co;
  FullAdder fa_s1_c14_r1(
    .io_a(fa_s1_c14_r1_io_a),
    .io_b(fa_s1_c14_r1_io_b),
    .io_ci(fa_s1_c14_r1_io_ci),
    .io_s(fa_s1_c14_r1_io_s),
    .io_co(fa_s1_c14_r1_io_co)
  );
  wire fa_s1_c14_r2_io_a;
  wire fa_s1_c14_r2_io_b;
  wire fa_s1_c14_r2_io_ci;
  wire fa_s1_c14_r2_io_s;
  wire fa_s1_c14_r2_io_co;
  FullAdder fa_s1_c14_r2(
    .io_a(fa_s1_c14_r2_io_a),
    .io_b(fa_s1_c14_r2_io_b),
    .io_ci(fa_s1_c14_r2_io_ci),
    .io_s(fa_s1_c14_r2_io_s),
    .io_co(fa_s1_c14_r2_io_co)
  );
  wire fa_s2_c14_r0_io_a;
  wire fa_s2_c14_r0_io_b;
  wire fa_s2_c14_r0_io_ci;
  wire fa_s2_c14_r0_io_s;
  wire fa_s2_c14_r0_io_co;
  FullAdder fa_s2_c14_r0(
    .io_a(fa_s2_c14_r0_io_a),
    .io_b(fa_s2_c14_r0_io_b),
    .io_ci(fa_s2_c14_r0_io_ci),
    .io_s(fa_s2_c14_r0_io_s),
    .io_co(fa_s2_c14_r0_io_co)
  );
  wire fa_s2_c14_r1_io_a;
  wire fa_s2_c14_r1_io_b;
  wire fa_s2_c14_r1_io_ci;
  wire fa_s2_c14_r1_io_s;
  wire fa_s2_c14_r1_io_co;
  FullAdder fa_s2_c14_r1(
    .io_a(fa_s2_c14_r1_io_a),
    .io_b(fa_s2_c14_r1_io_b),
    .io_ci(fa_s2_c14_r1_io_ci),
    .io_s(fa_s2_c14_r1_io_s),
    .io_co(fa_s2_c14_r1_io_co)
  );
  wire fa_s3_c14_r0_io_a;
  wire fa_s3_c14_r0_io_b;
  wire fa_s3_c14_r0_io_ci;
  wire fa_s3_c14_r0_io_s;
  wire fa_s3_c14_r0_io_co;
  FullAdder fa_s3_c14_r0(
    .io_a(fa_s3_c14_r0_io_a),
    .io_b(fa_s3_c14_r0_io_b),
    .io_ci(fa_s3_c14_r0_io_ci),
    .io_s(fa_s3_c14_r0_io_s),
    .io_co(fa_s3_c14_r0_io_co)
  );
  wire ft_s3_c14_r1_io_a;
  wire ft_s3_c14_r1_io_s;
  FallThrough ft_s3_c14_r1(
    .io_a(ft_s3_c14_r1_io_a),
    .io_s(ft_s3_c14_r1_io_s)
  );
  wire fa_s4_c14_r0_io_a;
  wire fa_s4_c14_r0_io_b;
  wire fa_s4_c14_r0_io_ci;
  wire fa_s4_c14_r0_io_s;
  wire fa_s4_c14_r0_io_co;
  FullAdder fa_s4_c14_r0(
    .io_a(fa_s4_c14_r0_io_a),
    .io_b(fa_s4_c14_r0_io_b),
    .io_ci(fa_s4_c14_r0_io_ci),
    .io_s(fa_s4_c14_r0_io_s),
    .io_co(fa_s4_c14_r0_io_co)
  );
  wire ft_s5_c14_r0_io_a;
  wire ft_s5_c14_r0_io_s;
  FallThrough ft_s5_c14_r0(
    .io_a(ft_s5_c14_r0_io_a),
    .io_s(ft_s5_c14_r0_io_s)
  );
  wire ft_s5_c14_r1_io_a;
  wire ft_s5_c14_r1_io_s;
  FallThrough ft_s5_c14_r1(
    .io_a(ft_s5_c14_r1_io_a),
    .io_s(ft_s5_c14_r1_io_s)
  );
  wire ft_s6_c14_r0_io_a;
  wire ft_s6_c14_r0_io_s;
  FallThrough ft_s6_c14_r0(
    .io_a(ft_s6_c14_r0_io_a),
    .io_s(ft_s6_c14_r0_io_s)
  );
  wire ft_s6_c14_r1_io_a;
  wire ft_s6_c14_r1_io_s;
  FallThrough ft_s6_c14_r1(
    .io_a(ft_s6_c14_r1_io_a),
    .io_s(ft_s6_c14_r1_io_s)
  );
  wire fa_s7_c14_r0_io_a;
  wire fa_s7_c14_r0_io_b;
  wire fa_s7_c14_r0_io_ci;
  wire fa_s7_c14_r0_io_s;
  wire fa_s7_c14_r0_io_co;
  FullAdder fa_s7_c14_r0(
    .io_a(fa_s7_c14_r0_io_a),
    .io_b(fa_s7_c14_r0_io_b),
    .io_ci(fa_s7_c14_r0_io_ci),
    .io_s(fa_s7_c14_r0_io_s),
    .io_co(fa_s7_c14_r0_io_co)
  );
  wire ft_s8_c14_r0_io_a;
  wire ft_s8_c14_r0_io_s;
  FallThrough ft_s8_c14_r0(
    .io_a(ft_s8_c14_r0_io_a),
    .io_s(ft_s8_c14_r0_io_s)
  );
  wire fa_s0_c15_r0_io_a;
  wire fa_s0_c15_r0_io_b;
  wire fa_s0_c15_r0_io_ci;
  wire fa_s0_c15_r0_io_s;
  wire fa_s0_c15_r0_io_co;
  FullAdder fa_s0_c15_r0(
    .io_a(fa_s0_c15_r0_io_a),
    .io_b(fa_s0_c15_r0_io_b),
    .io_ci(fa_s0_c15_r0_io_ci),
    .io_s(fa_s0_c15_r0_io_s),
    .io_co(fa_s0_c15_r0_io_co)
  );
  wire fa_s0_c15_r1_io_a;
  wire fa_s0_c15_r1_io_b;
  wire fa_s0_c15_r1_io_ci;
  wire fa_s0_c15_r1_io_s;
  wire fa_s0_c15_r1_io_co;
  FullAdder fa_s0_c15_r1(
    .io_a(fa_s0_c15_r1_io_a),
    .io_b(fa_s0_c15_r1_io_b),
    .io_ci(fa_s0_c15_r1_io_ci),
    .io_s(fa_s0_c15_r1_io_s),
    .io_co(fa_s0_c15_r1_io_co)
  );
  wire fa_s0_c15_r2_io_a;
  wire fa_s0_c15_r2_io_b;
  wire fa_s0_c15_r2_io_ci;
  wire fa_s0_c15_r2_io_s;
  wire fa_s0_c15_r2_io_co;
  FullAdder fa_s0_c15_r2(
    .io_a(fa_s0_c15_r2_io_a),
    .io_b(fa_s0_c15_r2_io_b),
    .io_ci(fa_s0_c15_r2_io_ci),
    .io_s(fa_s0_c15_r2_io_s),
    .io_co(fa_s0_c15_r2_io_co)
  );
  wire fa_s0_c15_r3_io_a;
  wire fa_s0_c15_r3_io_b;
  wire fa_s0_c15_r3_io_ci;
  wire fa_s0_c15_r3_io_s;
  wire fa_s0_c15_r3_io_co;
  FullAdder fa_s0_c15_r3(
    .io_a(fa_s0_c15_r3_io_a),
    .io_b(fa_s0_c15_r3_io_b),
    .io_ci(fa_s0_c15_r3_io_ci),
    .io_s(fa_s0_c15_r3_io_s),
    .io_co(fa_s0_c15_r3_io_co)
  );
  wire fa_s0_c15_r4_io_a;
  wire fa_s0_c15_r4_io_b;
  wire fa_s0_c15_r4_io_ci;
  wire fa_s0_c15_r4_io_s;
  wire fa_s0_c15_r4_io_co;
  FullAdder fa_s0_c15_r4(
    .io_a(fa_s0_c15_r4_io_a),
    .io_b(fa_s0_c15_r4_io_b),
    .io_ci(fa_s0_c15_r4_io_ci),
    .io_s(fa_s0_c15_r4_io_s),
    .io_co(fa_s0_c15_r4_io_co)
  );
  wire ft_s0_c15_r5_io_a;
  wire ft_s0_c15_r5_io_s;
  FallThrough ft_s0_c15_r5(
    .io_a(ft_s0_c15_r5_io_a),
    .io_s(ft_s0_c15_r5_io_s)
  );
  wire fa_s1_c15_r0_io_a;
  wire fa_s1_c15_r0_io_b;
  wire fa_s1_c15_r0_io_ci;
  wire fa_s1_c15_r0_io_s;
  wire fa_s1_c15_r0_io_co;
  FullAdder fa_s1_c15_r0(
    .io_a(fa_s1_c15_r0_io_a),
    .io_b(fa_s1_c15_r0_io_b),
    .io_ci(fa_s1_c15_r0_io_ci),
    .io_s(fa_s1_c15_r0_io_s),
    .io_co(fa_s1_c15_r0_io_co)
  );
  wire fa_s1_c15_r1_io_a;
  wire fa_s1_c15_r1_io_b;
  wire fa_s1_c15_r1_io_ci;
  wire fa_s1_c15_r1_io_s;
  wire fa_s1_c15_r1_io_co;
  FullAdder fa_s1_c15_r1(
    .io_a(fa_s1_c15_r1_io_a),
    .io_b(fa_s1_c15_r1_io_b),
    .io_ci(fa_s1_c15_r1_io_ci),
    .io_s(fa_s1_c15_r1_io_s),
    .io_co(fa_s1_c15_r1_io_co)
  );
  wire fa_s1_c15_r2_io_a;
  wire fa_s1_c15_r2_io_b;
  wire fa_s1_c15_r2_io_ci;
  wire fa_s1_c15_r2_io_s;
  wire fa_s1_c15_r2_io_co;
  FullAdder fa_s1_c15_r2(
    .io_a(fa_s1_c15_r2_io_a),
    .io_b(fa_s1_c15_r2_io_b),
    .io_ci(fa_s1_c15_r2_io_ci),
    .io_s(fa_s1_c15_r2_io_s),
    .io_co(fa_s1_c15_r2_io_co)
  );
  wire ha_s1_c15_r3_io_a;
  wire ha_s1_c15_r3_io_b;
  wire ha_s1_c15_r3_io_s;
  wire ha_s1_c15_r3_io_co;
  HalfAdder ha_s1_c15_r3(
    .io_a(ha_s1_c15_r3_io_a),
    .io_b(ha_s1_c15_r3_io_b),
    .io_s(ha_s1_c15_r3_io_s),
    .io_co(ha_s1_c15_r3_io_co)
  );
  wire fa_s2_c15_r0_io_a;
  wire fa_s2_c15_r0_io_b;
  wire fa_s2_c15_r0_io_ci;
  wire fa_s2_c15_r0_io_s;
  wire fa_s2_c15_r0_io_co;
  FullAdder fa_s2_c15_r0(
    .io_a(fa_s2_c15_r0_io_a),
    .io_b(fa_s2_c15_r0_io_b),
    .io_ci(fa_s2_c15_r0_io_ci),
    .io_s(fa_s2_c15_r0_io_s),
    .io_co(fa_s2_c15_r0_io_co)
  );
  wire fa_s2_c15_r1_io_a;
  wire fa_s2_c15_r1_io_b;
  wire fa_s2_c15_r1_io_ci;
  wire fa_s2_c15_r1_io_s;
  wire fa_s2_c15_r1_io_co;
  FullAdder fa_s2_c15_r1(
    .io_a(fa_s2_c15_r1_io_a),
    .io_b(fa_s2_c15_r1_io_b),
    .io_ci(fa_s2_c15_r1_io_ci),
    .io_s(fa_s2_c15_r1_io_s),
    .io_co(fa_s2_c15_r1_io_co)
  );
  wire ft_s2_c15_r2_io_a;
  wire ft_s2_c15_r2_io_s;
  FallThrough ft_s2_c15_r2(
    .io_a(ft_s2_c15_r2_io_a),
    .io_s(ft_s2_c15_r2_io_s)
  );
  wire fa_s3_c15_r0_io_a;
  wire fa_s3_c15_r0_io_b;
  wire fa_s3_c15_r0_io_ci;
  wire fa_s3_c15_r0_io_s;
  wire fa_s3_c15_r0_io_co;
  FullAdder fa_s3_c15_r0(
    .io_a(fa_s3_c15_r0_io_a),
    .io_b(fa_s3_c15_r0_io_b),
    .io_ci(fa_s3_c15_r0_io_ci),
    .io_s(fa_s3_c15_r0_io_s),
    .io_co(fa_s3_c15_r0_io_co)
  );
  wire ft_s3_c15_r1_io_a;
  wire ft_s3_c15_r1_io_s;
  FallThrough ft_s3_c15_r1(
    .io_a(ft_s3_c15_r1_io_a),
    .io_s(ft_s3_c15_r1_io_s)
  );
  wire ft_s3_c15_r2_io_a;
  wire ft_s3_c15_r2_io_s;
  FallThrough ft_s3_c15_r2(
    .io_a(ft_s3_c15_r2_io_a),
    .io_s(ft_s3_c15_r2_io_s)
  );
  wire fa_s4_c15_r0_io_a;
  wire fa_s4_c15_r0_io_b;
  wire fa_s4_c15_r0_io_ci;
  wire fa_s4_c15_r0_io_s;
  wire fa_s4_c15_r0_io_co;
  FullAdder fa_s4_c15_r0(
    .io_a(fa_s4_c15_r0_io_a),
    .io_b(fa_s4_c15_r0_io_b),
    .io_ci(fa_s4_c15_r0_io_ci),
    .io_s(fa_s4_c15_r0_io_s),
    .io_co(fa_s4_c15_r0_io_co)
  );
  wire ft_s4_c15_r1_io_a;
  wire ft_s4_c15_r1_io_s;
  FallThrough ft_s4_c15_r1(
    .io_a(ft_s4_c15_r1_io_a),
    .io_s(ft_s4_c15_r1_io_s)
  );
  wire fa_s5_c15_r0_io_a;
  wire fa_s5_c15_r0_io_b;
  wire fa_s5_c15_r0_io_ci;
  wire fa_s5_c15_r0_io_s;
  wire fa_s5_c15_r0_io_co;
  FullAdder fa_s5_c15_r0(
    .io_a(fa_s5_c15_r0_io_a),
    .io_b(fa_s5_c15_r0_io_b),
    .io_ci(fa_s5_c15_r0_io_ci),
    .io_s(fa_s5_c15_r0_io_s),
    .io_co(fa_s5_c15_r0_io_co)
  );
  wire ft_s6_c15_r0_io_a;
  wire ft_s6_c15_r0_io_s;
  FallThrough ft_s6_c15_r0(
    .io_a(ft_s6_c15_r0_io_a),
    .io_s(ft_s6_c15_r0_io_s)
  );
  wire ft_s7_c15_r0_io_a;
  wire ft_s7_c15_r0_io_s;
  FallThrough ft_s7_c15_r0(
    .io_a(ft_s7_c15_r0_io_a),
    .io_s(ft_s7_c15_r0_io_s)
  );
  wire ft_s8_c15_r0_io_a;
  wire ft_s8_c15_r0_io_s;
  FallThrough ft_s8_c15_r0(
    .io_a(ft_s8_c15_r0_io_a),
    .io_s(ft_s8_c15_r0_io_s)
  );
  wire ft_s8_c15_r1_io_a;
  wire ft_s8_c15_r1_io_s;
  FallThrough ft_s8_c15_r1(
    .io_a(ft_s8_c15_r1_io_a),
    .io_s(ft_s8_c15_r1_io_s)
  );
  wire fa_s0_c16_r0_io_a;
  wire fa_s0_c16_r0_io_b;
  wire fa_s0_c16_r0_io_ci;
  wire fa_s0_c16_r0_io_s;
  wire fa_s0_c16_r0_io_co;
  FullAdder fa_s0_c16_r0(
    .io_a(fa_s0_c16_r0_io_a),
    .io_b(fa_s0_c16_r0_io_b),
    .io_ci(fa_s0_c16_r0_io_ci),
    .io_s(fa_s0_c16_r0_io_s),
    .io_co(fa_s0_c16_r0_io_co)
  );
  wire fa_s0_c16_r1_io_a;
  wire fa_s0_c16_r1_io_b;
  wire fa_s0_c16_r1_io_ci;
  wire fa_s0_c16_r1_io_s;
  wire fa_s0_c16_r1_io_co;
  FullAdder fa_s0_c16_r1(
    .io_a(fa_s0_c16_r1_io_a),
    .io_b(fa_s0_c16_r1_io_b),
    .io_ci(fa_s0_c16_r1_io_ci),
    .io_s(fa_s0_c16_r1_io_s),
    .io_co(fa_s0_c16_r1_io_co)
  );
  wire fa_s0_c16_r2_io_a;
  wire fa_s0_c16_r2_io_b;
  wire fa_s0_c16_r2_io_ci;
  wire fa_s0_c16_r2_io_s;
  wire fa_s0_c16_r2_io_co;
  FullAdder fa_s0_c16_r2(
    .io_a(fa_s0_c16_r2_io_a),
    .io_b(fa_s0_c16_r2_io_b),
    .io_ci(fa_s0_c16_r2_io_ci),
    .io_s(fa_s0_c16_r2_io_s),
    .io_co(fa_s0_c16_r2_io_co)
  );
  wire fa_s0_c16_r3_io_a;
  wire fa_s0_c16_r3_io_b;
  wire fa_s0_c16_r3_io_ci;
  wire fa_s0_c16_r3_io_s;
  wire fa_s0_c16_r3_io_co;
  FullAdder fa_s0_c16_r3(
    .io_a(fa_s0_c16_r3_io_a),
    .io_b(fa_s0_c16_r3_io_b),
    .io_ci(fa_s0_c16_r3_io_ci),
    .io_s(fa_s0_c16_r3_io_s),
    .io_co(fa_s0_c16_r3_io_co)
  );
  wire fa_s0_c16_r4_io_a;
  wire fa_s0_c16_r4_io_b;
  wire fa_s0_c16_r4_io_ci;
  wire fa_s0_c16_r4_io_s;
  wire fa_s0_c16_r4_io_co;
  FullAdder fa_s0_c16_r4(
    .io_a(fa_s0_c16_r4_io_a),
    .io_b(fa_s0_c16_r4_io_b),
    .io_ci(fa_s0_c16_r4_io_ci),
    .io_s(fa_s0_c16_r4_io_s),
    .io_co(fa_s0_c16_r4_io_co)
  );
  wire fa_s1_c16_r0_io_a;
  wire fa_s1_c16_r0_io_b;
  wire fa_s1_c16_r0_io_ci;
  wire fa_s1_c16_r0_io_s;
  wire fa_s1_c16_r0_io_co;
  FullAdder fa_s1_c16_r0(
    .io_a(fa_s1_c16_r0_io_a),
    .io_b(fa_s1_c16_r0_io_b),
    .io_ci(fa_s1_c16_r0_io_ci),
    .io_s(fa_s1_c16_r0_io_s),
    .io_co(fa_s1_c16_r0_io_co)
  );
  wire fa_s1_c16_r1_io_a;
  wire fa_s1_c16_r1_io_b;
  wire fa_s1_c16_r1_io_ci;
  wire fa_s1_c16_r1_io_s;
  wire fa_s1_c16_r1_io_co;
  FullAdder fa_s1_c16_r1(
    .io_a(fa_s1_c16_r1_io_a),
    .io_b(fa_s1_c16_r1_io_b),
    .io_ci(fa_s1_c16_r1_io_ci),
    .io_s(fa_s1_c16_r1_io_s),
    .io_co(fa_s1_c16_r1_io_co)
  );
  wire fa_s1_c16_r2_io_a;
  wire fa_s1_c16_r2_io_b;
  wire fa_s1_c16_r2_io_ci;
  wire fa_s1_c16_r2_io_s;
  wire fa_s1_c16_r2_io_co;
  FullAdder fa_s1_c16_r2(
    .io_a(fa_s1_c16_r2_io_a),
    .io_b(fa_s1_c16_r2_io_b),
    .io_ci(fa_s1_c16_r2_io_ci),
    .io_s(fa_s1_c16_r2_io_s),
    .io_co(fa_s1_c16_r2_io_co)
  );
  wire ft_s1_c16_r3_io_a;
  wire ft_s1_c16_r3_io_s;
  FallThrough ft_s1_c16_r3(
    .io_a(ft_s1_c16_r3_io_a),
    .io_s(ft_s1_c16_r3_io_s)
  );
  wire fa_s2_c16_r0_io_a;
  wire fa_s2_c16_r0_io_b;
  wire fa_s2_c16_r0_io_ci;
  wire fa_s2_c16_r0_io_s;
  wire fa_s2_c16_r0_io_co;
  FullAdder fa_s2_c16_r0(
    .io_a(fa_s2_c16_r0_io_a),
    .io_b(fa_s2_c16_r0_io_b),
    .io_ci(fa_s2_c16_r0_io_ci),
    .io_s(fa_s2_c16_r0_io_s),
    .io_co(fa_s2_c16_r0_io_co)
  );
  wire fa_s2_c16_r1_io_a;
  wire fa_s2_c16_r1_io_b;
  wire fa_s2_c16_r1_io_ci;
  wire fa_s2_c16_r1_io_s;
  wire fa_s2_c16_r1_io_co;
  FullAdder fa_s2_c16_r1(
    .io_a(fa_s2_c16_r1_io_a),
    .io_b(fa_s2_c16_r1_io_b),
    .io_ci(fa_s2_c16_r1_io_ci),
    .io_s(fa_s2_c16_r1_io_s),
    .io_co(fa_s2_c16_r1_io_co)
  );
  wire ha_s2_c16_r2_io_a;
  wire ha_s2_c16_r2_io_b;
  wire ha_s2_c16_r2_io_s;
  wire ha_s2_c16_r2_io_co;
  HalfAdder ha_s2_c16_r2(
    .io_a(ha_s2_c16_r2_io_a),
    .io_b(ha_s2_c16_r2_io_b),
    .io_s(ha_s2_c16_r2_io_s),
    .io_co(ha_s2_c16_r2_io_co)
  );
  wire fa_s3_c16_r0_io_a;
  wire fa_s3_c16_r0_io_b;
  wire fa_s3_c16_r0_io_ci;
  wire fa_s3_c16_r0_io_s;
  wire fa_s3_c16_r0_io_co;
  FullAdder fa_s3_c16_r0(
    .io_a(fa_s3_c16_r0_io_a),
    .io_b(fa_s3_c16_r0_io_b),
    .io_ci(fa_s3_c16_r0_io_ci),
    .io_s(fa_s3_c16_r0_io_s),
    .io_co(fa_s3_c16_r0_io_co)
  );
  wire ft_s3_c16_r1_io_a;
  wire ft_s3_c16_r1_io_s;
  FallThrough ft_s3_c16_r1(
    .io_a(ft_s3_c16_r1_io_a),
    .io_s(ft_s3_c16_r1_io_s)
  );
  wire ft_s3_c16_r2_io_a;
  wire ft_s3_c16_r2_io_s;
  FallThrough ft_s3_c16_r2(
    .io_a(ft_s3_c16_r2_io_a),
    .io_s(ft_s3_c16_r2_io_s)
  );
  wire fa_s4_c16_r0_io_a;
  wire fa_s4_c16_r0_io_b;
  wire fa_s4_c16_r0_io_ci;
  wire fa_s4_c16_r0_io_s;
  wire fa_s4_c16_r0_io_co;
  FullAdder fa_s4_c16_r0(
    .io_a(fa_s4_c16_r0_io_a),
    .io_b(fa_s4_c16_r0_io_b),
    .io_ci(fa_s4_c16_r0_io_ci),
    .io_s(fa_s4_c16_r0_io_s),
    .io_co(fa_s4_c16_r0_io_co)
  );
  wire ft_s4_c16_r1_io_a;
  wire ft_s4_c16_r1_io_s;
  FallThrough ft_s4_c16_r1(
    .io_a(ft_s4_c16_r1_io_a),
    .io_s(ft_s4_c16_r1_io_s)
  );
  wire fa_s5_c16_r0_io_a;
  wire fa_s5_c16_r0_io_b;
  wire fa_s5_c16_r0_io_ci;
  wire fa_s5_c16_r0_io_s;
  wire fa_s5_c16_r0_io_co;
  FullAdder fa_s5_c16_r0(
    .io_a(fa_s5_c16_r0_io_a),
    .io_b(fa_s5_c16_r0_io_b),
    .io_ci(fa_s5_c16_r0_io_ci),
    .io_s(fa_s5_c16_r0_io_s),
    .io_co(fa_s5_c16_r0_io_co)
  );
  wire ft_s6_c16_r0_io_a;
  wire ft_s6_c16_r0_io_s;
  FallThrough ft_s6_c16_r0(
    .io_a(ft_s6_c16_r0_io_a),
    .io_s(ft_s6_c16_r0_io_s)
  );
  wire ft_s6_c16_r1_io_a;
  wire ft_s6_c16_r1_io_s;
  FallThrough ft_s6_c16_r1(
    .io_a(ft_s6_c16_r1_io_a),
    .io_s(ft_s6_c16_r1_io_s)
  );
  wire ft_s7_c16_r0_io_a;
  wire ft_s7_c16_r0_io_s;
  FallThrough ft_s7_c16_r0(
    .io_a(ft_s7_c16_r0_io_a),
    .io_s(ft_s7_c16_r0_io_s)
  );
  wire ft_s7_c16_r1_io_a;
  wire ft_s7_c16_r1_io_s;
  FallThrough ft_s7_c16_r1(
    .io_a(ft_s7_c16_r1_io_a),
    .io_s(ft_s7_c16_r1_io_s)
  );
  wire ft_s8_c16_r0_io_a;
  wire ft_s8_c16_r0_io_s;
  FallThrough ft_s8_c16_r0(
    .io_a(ft_s8_c16_r0_io_a),
    .io_s(ft_s8_c16_r0_io_s)
  );
  wire ft_s8_c16_r1_io_a;
  wire ft_s8_c16_r1_io_s;
  FallThrough ft_s8_c16_r1(
    .io_a(ft_s8_c16_r1_io_a),
    .io_s(ft_s8_c16_r1_io_s)
  );
  wire fa_s0_c17_r0_io_a;
  wire fa_s0_c17_r0_io_b;
  wire fa_s0_c17_r0_io_ci;
  wire fa_s0_c17_r0_io_s;
  wire fa_s0_c17_r0_io_co;
  FullAdder fa_s0_c17_r0(
    .io_a(fa_s0_c17_r0_io_a),
    .io_b(fa_s0_c17_r0_io_b),
    .io_ci(fa_s0_c17_r0_io_ci),
    .io_s(fa_s0_c17_r0_io_s),
    .io_co(fa_s0_c17_r0_io_co)
  );
  wire fa_s0_c17_r1_io_a;
  wire fa_s0_c17_r1_io_b;
  wire fa_s0_c17_r1_io_ci;
  wire fa_s0_c17_r1_io_s;
  wire fa_s0_c17_r1_io_co;
  FullAdder fa_s0_c17_r1(
    .io_a(fa_s0_c17_r1_io_a),
    .io_b(fa_s0_c17_r1_io_b),
    .io_ci(fa_s0_c17_r1_io_ci),
    .io_s(fa_s0_c17_r1_io_s),
    .io_co(fa_s0_c17_r1_io_co)
  );
  wire fa_s0_c17_r2_io_a;
  wire fa_s0_c17_r2_io_b;
  wire fa_s0_c17_r2_io_ci;
  wire fa_s0_c17_r2_io_s;
  wire fa_s0_c17_r2_io_co;
  FullAdder fa_s0_c17_r2(
    .io_a(fa_s0_c17_r2_io_a),
    .io_b(fa_s0_c17_r2_io_b),
    .io_ci(fa_s0_c17_r2_io_ci),
    .io_s(fa_s0_c17_r2_io_s),
    .io_co(fa_s0_c17_r2_io_co)
  );
  wire fa_s0_c17_r3_io_a;
  wire fa_s0_c17_r3_io_b;
  wire fa_s0_c17_r3_io_ci;
  wire fa_s0_c17_r3_io_s;
  wire fa_s0_c17_r3_io_co;
  FullAdder fa_s0_c17_r3(
    .io_a(fa_s0_c17_r3_io_a),
    .io_b(fa_s0_c17_r3_io_b),
    .io_ci(fa_s0_c17_r3_io_ci),
    .io_s(fa_s0_c17_r3_io_s),
    .io_co(fa_s0_c17_r3_io_co)
  );
  wire ft_s0_c17_r4_io_a;
  wire ft_s0_c17_r4_io_s;
  FallThrough ft_s0_c17_r4(
    .io_a(ft_s0_c17_r4_io_a),
    .io_s(ft_s0_c17_r4_io_s)
  );
  wire ft_s0_c17_r5_io_a;
  wire ft_s0_c17_r5_io_s;
  FallThrough ft_s0_c17_r5(
    .io_a(ft_s0_c17_r5_io_a),
    .io_s(ft_s0_c17_r5_io_s)
  );
  wire fa_s1_c17_r0_io_a;
  wire fa_s1_c17_r0_io_b;
  wire fa_s1_c17_r0_io_ci;
  wire fa_s1_c17_r0_io_s;
  wire fa_s1_c17_r0_io_co;
  FullAdder fa_s1_c17_r0(
    .io_a(fa_s1_c17_r0_io_a),
    .io_b(fa_s1_c17_r0_io_b),
    .io_ci(fa_s1_c17_r0_io_ci),
    .io_s(fa_s1_c17_r0_io_s),
    .io_co(fa_s1_c17_r0_io_co)
  );
  wire fa_s1_c17_r1_io_a;
  wire fa_s1_c17_r1_io_b;
  wire fa_s1_c17_r1_io_ci;
  wire fa_s1_c17_r1_io_s;
  wire fa_s1_c17_r1_io_co;
  FullAdder fa_s1_c17_r1(
    .io_a(fa_s1_c17_r1_io_a),
    .io_b(fa_s1_c17_r1_io_b),
    .io_ci(fa_s1_c17_r1_io_ci),
    .io_s(fa_s1_c17_r1_io_s),
    .io_co(fa_s1_c17_r1_io_co)
  );
  wire fa_s1_c17_r2_io_a;
  wire fa_s1_c17_r2_io_b;
  wire fa_s1_c17_r2_io_ci;
  wire fa_s1_c17_r2_io_s;
  wire fa_s1_c17_r2_io_co;
  FullAdder fa_s1_c17_r2(
    .io_a(fa_s1_c17_r2_io_a),
    .io_b(fa_s1_c17_r2_io_b),
    .io_ci(fa_s1_c17_r2_io_ci),
    .io_s(fa_s1_c17_r2_io_s),
    .io_co(fa_s1_c17_r2_io_co)
  );
  wire ft_s1_c17_r3_io_a;
  wire ft_s1_c17_r3_io_s;
  FallThrough ft_s1_c17_r3(
    .io_a(ft_s1_c17_r3_io_a),
    .io_s(ft_s1_c17_r3_io_s)
  );
  wire ft_s1_c17_r4_io_a;
  wire ft_s1_c17_r4_io_s;
  FallThrough ft_s1_c17_r4(
    .io_a(ft_s1_c17_r4_io_a),
    .io_s(ft_s1_c17_r4_io_s)
  );
  wire fa_s2_c17_r0_io_a;
  wire fa_s2_c17_r0_io_b;
  wire fa_s2_c17_r0_io_ci;
  wire fa_s2_c17_r0_io_s;
  wire fa_s2_c17_r0_io_co;
  FullAdder fa_s2_c17_r0(
    .io_a(fa_s2_c17_r0_io_a),
    .io_b(fa_s2_c17_r0_io_b),
    .io_ci(fa_s2_c17_r0_io_ci),
    .io_s(fa_s2_c17_r0_io_s),
    .io_co(fa_s2_c17_r0_io_co)
  );
  wire fa_s2_c17_r1_io_a;
  wire fa_s2_c17_r1_io_b;
  wire fa_s2_c17_r1_io_ci;
  wire fa_s2_c17_r1_io_s;
  wire fa_s2_c17_r1_io_co;
  FullAdder fa_s2_c17_r1(
    .io_a(fa_s2_c17_r1_io_a),
    .io_b(fa_s2_c17_r1_io_b),
    .io_ci(fa_s2_c17_r1_io_ci),
    .io_s(fa_s2_c17_r1_io_s),
    .io_co(fa_s2_c17_r1_io_co)
  );
  wire ft_s2_c17_r2_io_a;
  wire ft_s2_c17_r2_io_s;
  FallThrough ft_s2_c17_r2(
    .io_a(ft_s2_c17_r2_io_a),
    .io_s(ft_s2_c17_r2_io_s)
  );
  wire ft_s2_c17_r3_io_a;
  wire ft_s2_c17_r3_io_s;
  FallThrough ft_s2_c17_r3(
    .io_a(ft_s2_c17_r3_io_a),
    .io_s(ft_s2_c17_r3_io_s)
  );
  wire fa_s3_c17_r0_io_a;
  wire fa_s3_c17_r0_io_b;
  wire fa_s3_c17_r0_io_ci;
  wire fa_s3_c17_r0_io_s;
  wire fa_s3_c17_r0_io_co;
  FullAdder fa_s3_c17_r0(
    .io_a(fa_s3_c17_r0_io_a),
    .io_b(fa_s3_c17_r0_io_b),
    .io_ci(fa_s3_c17_r0_io_ci),
    .io_s(fa_s3_c17_r0_io_s),
    .io_co(fa_s3_c17_r0_io_co)
  );
  wire fa_s3_c17_r1_io_a;
  wire fa_s3_c17_r1_io_b;
  wire fa_s3_c17_r1_io_ci;
  wire fa_s3_c17_r1_io_s;
  wire fa_s3_c17_r1_io_co;
  FullAdder fa_s3_c17_r1(
    .io_a(fa_s3_c17_r1_io_a),
    .io_b(fa_s3_c17_r1_io_b),
    .io_ci(fa_s3_c17_r1_io_ci),
    .io_s(fa_s3_c17_r1_io_s),
    .io_co(fa_s3_c17_r1_io_co)
  );
  wire ft_s3_c17_r2_io_a;
  wire ft_s3_c17_r2_io_s;
  FallThrough ft_s3_c17_r2(
    .io_a(ft_s3_c17_r2_io_a),
    .io_s(ft_s3_c17_r2_io_s)
  );
  wire fa_s4_c17_r0_io_a;
  wire fa_s4_c17_r0_io_b;
  wire fa_s4_c17_r0_io_ci;
  wire fa_s4_c17_r0_io_s;
  wire fa_s4_c17_r0_io_co;
  FullAdder fa_s4_c17_r0(
    .io_a(fa_s4_c17_r0_io_a),
    .io_b(fa_s4_c17_r0_io_b),
    .io_ci(fa_s4_c17_r0_io_ci),
    .io_s(fa_s4_c17_r0_io_s),
    .io_co(fa_s4_c17_r0_io_co)
  );
  wire ft_s4_c17_r1_io_a;
  wire ft_s4_c17_r1_io_s;
  FallThrough ft_s4_c17_r1(
    .io_a(ft_s4_c17_r1_io_a),
    .io_s(ft_s4_c17_r1_io_s)
  );
  wire fa_s5_c17_r0_io_a;
  wire fa_s5_c17_r0_io_b;
  wire fa_s5_c17_r0_io_ci;
  wire fa_s5_c17_r0_io_s;
  wire fa_s5_c17_r0_io_co;
  FullAdder fa_s5_c17_r0(
    .io_a(fa_s5_c17_r0_io_a),
    .io_b(fa_s5_c17_r0_io_b),
    .io_ci(fa_s5_c17_r0_io_ci),
    .io_s(fa_s5_c17_r0_io_s),
    .io_co(fa_s5_c17_r0_io_co)
  );
  wire ft_s6_c17_r0_io_a;
  wire ft_s6_c17_r0_io_s;
  FallThrough ft_s6_c17_r0(
    .io_a(ft_s6_c17_r0_io_a),
    .io_s(ft_s6_c17_r0_io_s)
  );
  wire ft_s6_c17_r1_io_a;
  wire ft_s6_c17_r1_io_s;
  FallThrough ft_s6_c17_r1(
    .io_a(ft_s6_c17_r1_io_a),
    .io_s(ft_s6_c17_r1_io_s)
  );
  wire ft_s7_c17_r0_io_a;
  wire ft_s7_c17_r0_io_s;
  FallThrough ft_s7_c17_r0(
    .io_a(ft_s7_c17_r0_io_a),
    .io_s(ft_s7_c17_r0_io_s)
  );
  wire ft_s7_c17_r1_io_a;
  wire ft_s7_c17_r1_io_s;
  FallThrough ft_s7_c17_r1(
    .io_a(ft_s7_c17_r1_io_a),
    .io_s(ft_s7_c17_r1_io_s)
  );
  wire ft_s8_c17_r0_io_a;
  wire ft_s8_c17_r0_io_s;
  FallThrough ft_s8_c17_r0(
    .io_a(ft_s8_c17_r0_io_a),
    .io_s(ft_s8_c17_r0_io_s)
  );
  wire ft_s8_c17_r1_io_a;
  wire ft_s8_c17_r1_io_s;
  FallThrough ft_s8_c17_r1(
    .io_a(ft_s8_c17_r1_io_a),
    .io_s(ft_s8_c17_r1_io_s)
  );
  wire fa_s0_c18_r0_io_a;
  wire fa_s0_c18_r0_io_b;
  wire fa_s0_c18_r0_io_ci;
  wire fa_s0_c18_r0_io_s;
  wire fa_s0_c18_r0_io_co;
  FullAdder fa_s0_c18_r0(
    .io_a(fa_s0_c18_r0_io_a),
    .io_b(fa_s0_c18_r0_io_b),
    .io_ci(fa_s0_c18_r0_io_ci),
    .io_s(fa_s0_c18_r0_io_s),
    .io_co(fa_s0_c18_r0_io_co)
  );
  wire fa_s0_c18_r1_io_a;
  wire fa_s0_c18_r1_io_b;
  wire fa_s0_c18_r1_io_ci;
  wire fa_s0_c18_r1_io_s;
  wire fa_s0_c18_r1_io_co;
  FullAdder fa_s0_c18_r1(
    .io_a(fa_s0_c18_r1_io_a),
    .io_b(fa_s0_c18_r1_io_b),
    .io_ci(fa_s0_c18_r1_io_ci),
    .io_s(fa_s0_c18_r1_io_s),
    .io_co(fa_s0_c18_r1_io_co)
  );
  wire fa_s0_c18_r2_io_a;
  wire fa_s0_c18_r2_io_b;
  wire fa_s0_c18_r2_io_ci;
  wire fa_s0_c18_r2_io_s;
  wire fa_s0_c18_r2_io_co;
  FullAdder fa_s0_c18_r2(
    .io_a(fa_s0_c18_r2_io_a),
    .io_b(fa_s0_c18_r2_io_b),
    .io_ci(fa_s0_c18_r2_io_ci),
    .io_s(fa_s0_c18_r2_io_s),
    .io_co(fa_s0_c18_r2_io_co)
  );
  wire fa_s0_c18_r3_io_a;
  wire fa_s0_c18_r3_io_b;
  wire fa_s0_c18_r3_io_ci;
  wire fa_s0_c18_r3_io_s;
  wire fa_s0_c18_r3_io_co;
  FullAdder fa_s0_c18_r3(
    .io_a(fa_s0_c18_r3_io_a),
    .io_b(fa_s0_c18_r3_io_b),
    .io_ci(fa_s0_c18_r3_io_ci),
    .io_s(fa_s0_c18_r3_io_s),
    .io_co(fa_s0_c18_r3_io_co)
  );
  wire ft_s0_c18_r4_io_a;
  wire ft_s0_c18_r4_io_s;
  FallThrough ft_s0_c18_r4(
    .io_a(ft_s0_c18_r4_io_a),
    .io_s(ft_s0_c18_r4_io_s)
  );
  wire fa_s1_c18_r0_io_a;
  wire fa_s1_c18_r0_io_b;
  wire fa_s1_c18_r0_io_ci;
  wire fa_s1_c18_r0_io_s;
  wire fa_s1_c18_r0_io_co;
  FullAdder fa_s1_c18_r0(
    .io_a(fa_s1_c18_r0_io_a),
    .io_b(fa_s1_c18_r0_io_b),
    .io_ci(fa_s1_c18_r0_io_ci),
    .io_s(fa_s1_c18_r0_io_s),
    .io_co(fa_s1_c18_r0_io_co)
  );
  wire fa_s1_c18_r1_io_a;
  wire fa_s1_c18_r1_io_b;
  wire fa_s1_c18_r1_io_ci;
  wire fa_s1_c18_r1_io_s;
  wire fa_s1_c18_r1_io_co;
  FullAdder fa_s1_c18_r1(
    .io_a(fa_s1_c18_r1_io_a),
    .io_b(fa_s1_c18_r1_io_b),
    .io_ci(fa_s1_c18_r1_io_ci),
    .io_s(fa_s1_c18_r1_io_s),
    .io_co(fa_s1_c18_r1_io_co)
  );
  wire fa_s1_c18_r2_io_a;
  wire fa_s1_c18_r2_io_b;
  wire fa_s1_c18_r2_io_ci;
  wire fa_s1_c18_r2_io_s;
  wire fa_s1_c18_r2_io_co;
  FullAdder fa_s1_c18_r2(
    .io_a(fa_s1_c18_r2_io_a),
    .io_b(fa_s1_c18_r2_io_b),
    .io_ci(fa_s1_c18_r2_io_ci),
    .io_s(fa_s1_c18_r2_io_s),
    .io_co(fa_s1_c18_r2_io_co)
  );
  wire fa_s2_c18_r0_io_a;
  wire fa_s2_c18_r0_io_b;
  wire fa_s2_c18_r0_io_ci;
  wire fa_s2_c18_r0_io_s;
  wire fa_s2_c18_r0_io_co;
  FullAdder fa_s2_c18_r0(
    .io_a(fa_s2_c18_r0_io_a),
    .io_b(fa_s2_c18_r0_io_b),
    .io_ci(fa_s2_c18_r0_io_ci),
    .io_s(fa_s2_c18_r0_io_s),
    .io_co(fa_s2_c18_r0_io_co)
  );
  wire fa_s2_c18_r1_io_a;
  wire fa_s2_c18_r1_io_b;
  wire fa_s2_c18_r1_io_ci;
  wire fa_s2_c18_r1_io_s;
  wire fa_s2_c18_r1_io_co;
  FullAdder fa_s2_c18_r1(
    .io_a(fa_s2_c18_r1_io_a),
    .io_b(fa_s2_c18_r1_io_b),
    .io_ci(fa_s2_c18_r1_io_ci),
    .io_s(fa_s2_c18_r1_io_s),
    .io_co(fa_s2_c18_r1_io_co)
  );
  wire fa_s3_c18_r0_io_a;
  wire fa_s3_c18_r0_io_b;
  wire fa_s3_c18_r0_io_ci;
  wire fa_s3_c18_r0_io_s;
  wire fa_s3_c18_r0_io_co;
  FullAdder fa_s3_c18_r0(
    .io_a(fa_s3_c18_r0_io_a),
    .io_b(fa_s3_c18_r0_io_b),
    .io_ci(fa_s3_c18_r0_io_ci),
    .io_s(fa_s3_c18_r0_io_s),
    .io_co(fa_s3_c18_r0_io_co)
  );
  wire ft_s3_c18_r1_io_a;
  wire ft_s3_c18_r1_io_s;
  FallThrough ft_s3_c18_r1(
    .io_a(ft_s3_c18_r1_io_a),
    .io_s(ft_s3_c18_r1_io_s)
  );
  wire fa_s4_c18_r0_io_a;
  wire fa_s4_c18_r0_io_b;
  wire fa_s4_c18_r0_io_ci;
  wire fa_s4_c18_r0_io_s;
  wire fa_s4_c18_r0_io_co;
  FullAdder fa_s4_c18_r0(
    .io_a(fa_s4_c18_r0_io_a),
    .io_b(fa_s4_c18_r0_io_b),
    .io_ci(fa_s4_c18_r0_io_ci),
    .io_s(fa_s4_c18_r0_io_s),
    .io_co(fa_s4_c18_r0_io_co)
  );
  wire ft_s4_c18_r1_io_a;
  wire ft_s4_c18_r1_io_s;
  FallThrough ft_s4_c18_r1(
    .io_a(ft_s4_c18_r1_io_a),
    .io_s(ft_s4_c18_r1_io_s)
  );
  wire fa_s5_c18_r0_io_a;
  wire fa_s5_c18_r0_io_b;
  wire fa_s5_c18_r0_io_ci;
  wire fa_s5_c18_r0_io_s;
  wire fa_s5_c18_r0_io_co;
  FullAdder fa_s5_c18_r0(
    .io_a(fa_s5_c18_r0_io_a),
    .io_b(fa_s5_c18_r0_io_b),
    .io_ci(fa_s5_c18_r0_io_ci),
    .io_s(fa_s5_c18_r0_io_s),
    .io_co(fa_s5_c18_r0_io_co)
  );
  wire ft_s6_c18_r0_io_a;
  wire ft_s6_c18_r0_io_s;
  FallThrough ft_s6_c18_r0(
    .io_a(ft_s6_c18_r0_io_a),
    .io_s(ft_s6_c18_r0_io_s)
  );
  wire ft_s6_c18_r1_io_a;
  wire ft_s6_c18_r1_io_s;
  FallThrough ft_s6_c18_r1(
    .io_a(ft_s6_c18_r1_io_a),
    .io_s(ft_s6_c18_r1_io_s)
  );
  wire ft_s7_c18_r0_io_a;
  wire ft_s7_c18_r0_io_s;
  FallThrough ft_s7_c18_r0(
    .io_a(ft_s7_c18_r0_io_a),
    .io_s(ft_s7_c18_r0_io_s)
  );
  wire ft_s7_c18_r1_io_a;
  wire ft_s7_c18_r1_io_s;
  FallThrough ft_s7_c18_r1(
    .io_a(ft_s7_c18_r1_io_a),
    .io_s(ft_s7_c18_r1_io_s)
  );
  wire ft_s8_c18_r0_io_a;
  wire ft_s8_c18_r0_io_s;
  FallThrough ft_s8_c18_r0(
    .io_a(ft_s8_c18_r0_io_a),
    .io_s(ft_s8_c18_r0_io_s)
  );
  wire ft_s8_c18_r1_io_a;
  wire ft_s8_c18_r1_io_s;
  FallThrough ft_s8_c18_r1(
    .io_a(ft_s8_c18_r1_io_a),
    .io_s(ft_s8_c18_r1_io_s)
  );
  wire fa_s0_c19_r0_io_a;
  wire fa_s0_c19_r0_io_b;
  wire fa_s0_c19_r0_io_ci;
  wire fa_s0_c19_r0_io_s;
  wire fa_s0_c19_r0_io_co;
  FullAdder fa_s0_c19_r0(
    .io_a(fa_s0_c19_r0_io_a),
    .io_b(fa_s0_c19_r0_io_b),
    .io_ci(fa_s0_c19_r0_io_ci),
    .io_s(fa_s0_c19_r0_io_s),
    .io_co(fa_s0_c19_r0_io_co)
  );
  wire fa_s0_c19_r1_io_a;
  wire fa_s0_c19_r1_io_b;
  wire fa_s0_c19_r1_io_ci;
  wire fa_s0_c19_r1_io_s;
  wire fa_s0_c19_r1_io_co;
  FullAdder fa_s0_c19_r1(
    .io_a(fa_s0_c19_r1_io_a),
    .io_b(fa_s0_c19_r1_io_b),
    .io_ci(fa_s0_c19_r1_io_ci),
    .io_s(fa_s0_c19_r1_io_s),
    .io_co(fa_s0_c19_r1_io_co)
  );
  wire fa_s0_c19_r2_io_a;
  wire fa_s0_c19_r2_io_b;
  wire fa_s0_c19_r2_io_ci;
  wire fa_s0_c19_r2_io_s;
  wire fa_s0_c19_r2_io_co;
  FullAdder fa_s0_c19_r2(
    .io_a(fa_s0_c19_r2_io_a),
    .io_b(fa_s0_c19_r2_io_b),
    .io_ci(fa_s0_c19_r2_io_ci),
    .io_s(fa_s0_c19_r2_io_s),
    .io_co(fa_s0_c19_r2_io_co)
  );
  wire fa_s0_c19_r3_io_a;
  wire fa_s0_c19_r3_io_b;
  wire fa_s0_c19_r3_io_ci;
  wire fa_s0_c19_r3_io_s;
  wire fa_s0_c19_r3_io_co;
  FullAdder fa_s0_c19_r3(
    .io_a(fa_s0_c19_r3_io_a),
    .io_b(fa_s0_c19_r3_io_b),
    .io_ci(fa_s0_c19_r3_io_ci),
    .io_s(fa_s0_c19_r3_io_s),
    .io_co(fa_s0_c19_r3_io_co)
  );
  wire fa_s1_c19_r0_io_a;
  wire fa_s1_c19_r0_io_b;
  wire fa_s1_c19_r0_io_ci;
  wire fa_s1_c19_r0_io_s;
  wire fa_s1_c19_r0_io_co;
  FullAdder fa_s1_c19_r0(
    .io_a(fa_s1_c19_r0_io_a),
    .io_b(fa_s1_c19_r0_io_b),
    .io_ci(fa_s1_c19_r0_io_ci),
    .io_s(fa_s1_c19_r0_io_s),
    .io_co(fa_s1_c19_r0_io_co)
  );
  wire fa_s1_c19_r1_io_a;
  wire fa_s1_c19_r1_io_b;
  wire fa_s1_c19_r1_io_ci;
  wire fa_s1_c19_r1_io_s;
  wire fa_s1_c19_r1_io_co;
  FullAdder fa_s1_c19_r1(
    .io_a(fa_s1_c19_r1_io_a),
    .io_b(fa_s1_c19_r1_io_b),
    .io_ci(fa_s1_c19_r1_io_ci),
    .io_s(fa_s1_c19_r1_io_s),
    .io_co(fa_s1_c19_r1_io_co)
  );
  wire ha_s1_c19_r2_io_a;
  wire ha_s1_c19_r2_io_b;
  wire ha_s1_c19_r2_io_s;
  wire ha_s1_c19_r2_io_co;
  HalfAdder ha_s1_c19_r2(
    .io_a(ha_s1_c19_r2_io_a),
    .io_b(ha_s1_c19_r2_io_b),
    .io_s(ha_s1_c19_r2_io_s),
    .io_co(ha_s1_c19_r2_io_co)
  );
  wire fa_s2_c19_r0_io_a;
  wire fa_s2_c19_r0_io_b;
  wire fa_s2_c19_r0_io_ci;
  wire fa_s2_c19_r0_io_s;
  wire fa_s2_c19_r0_io_co;
  FullAdder fa_s2_c19_r0(
    .io_a(fa_s2_c19_r0_io_a),
    .io_b(fa_s2_c19_r0_io_b),
    .io_ci(fa_s2_c19_r0_io_ci),
    .io_s(fa_s2_c19_r0_io_s),
    .io_co(fa_s2_c19_r0_io_co)
  );
  wire fa_s2_c19_r1_io_a;
  wire fa_s2_c19_r1_io_b;
  wire fa_s2_c19_r1_io_ci;
  wire fa_s2_c19_r1_io_s;
  wire fa_s2_c19_r1_io_co;
  FullAdder fa_s2_c19_r1(
    .io_a(fa_s2_c19_r1_io_a),
    .io_b(fa_s2_c19_r1_io_b),
    .io_ci(fa_s2_c19_r1_io_ci),
    .io_s(fa_s2_c19_r1_io_s),
    .io_co(fa_s2_c19_r1_io_co)
  );
  wire fa_s3_c19_r0_io_a;
  wire fa_s3_c19_r0_io_b;
  wire fa_s3_c19_r0_io_ci;
  wire fa_s3_c19_r0_io_s;
  wire fa_s3_c19_r0_io_co;
  FullAdder fa_s3_c19_r0(
    .io_a(fa_s3_c19_r0_io_a),
    .io_b(fa_s3_c19_r0_io_b),
    .io_ci(fa_s3_c19_r0_io_ci),
    .io_s(fa_s3_c19_r0_io_s),
    .io_co(fa_s3_c19_r0_io_co)
  );
  wire ft_s3_c19_r1_io_a;
  wire ft_s3_c19_r1_io_s;
  FallThrough ft_s3_c19_r1(
    .io_a(ft_s3_c19_r1_io_a),
    .io_s(ft_s3_c19_r1_io_s)
  );
  wire fa_s4_c19_r0_io_a;
  wire fa_s4_c19_r0_io_b;
  wire fa_s4_c19_r0_io_ci;
  wire fa_s4_c19_r0_io_s;
  wire fa_s4_c19_r0_io_co;
  FullAdder fa_s4_c19_r0(
    .io_a(fa_s4_c19_r0_io_a),
    .io_b(fa_s4_c19_r0_io_b),
    .io_ci(fa_s4_c19_r0_io_ci),
    .io_s(fa_s4_c19_r0_io_s),
    .io_co(fa_s4_c19_r0_io_co)
  );
  wire ft_s5_c19_r0_io_a;
  wire ft_s5_c19_r0_io_s;
  FallThrough ft_s5_c19_r0(
    .io_a(ft_s5_c19_r0_io_a),
    .io_s(ft_s5_c19_r0_io_s)
  );
  wire ft_s5_c19_r1_io_a;
  wire ft_s5_c19_r1_io_s;
  FallThrough ft_s5_c19_r1(
    .io_a(ft_s5_c19_r1_io_a),
    .io_s(ft_s5_c19_r1_io_s)
  );
  wire fa_s6_c19_r0_io_a;
  wire fa_s6_c19_r0_io_b;
  wire fa_s6_c19_r0_io_ci;
  wire fa_s6_c19_r0_io_s;
  wire fa_s6_c19_r0_io_co;
  FullAdder fa_s6_c19_r0(
    .io_a(fa_s6_c19_r0_io_a),
    .io_b(fa_s6_c19_r0_io_b),
    .io_ci(fa_s6_c19_r0_io_ci),
    .io_s(fa_s6_c19_r0_io_s),
    .io_co(fa_s6_c19_r0_io_co)
  );
  wire ft_s7_c19_r0_io_a;
  wire ft_s7_c19_r0_io_s;
  FallThrough ft_s7_c19_r0(
    .io_a(ft_s7_c19_r0_io_a),
    .io_s(ft_s7_c19_r0_io_s)
  );
  wire ft_s8_c19_r0_io_a;
  wire ft_s8_c19_r0_io_s;
  FallThrough ft_s8_c19_r0(
    .io_a(ft_s8_c19_r0_io_a),
    .io_s(ft_s8_c19_r0_io_s)
  );
  wire fa_s0_c20_r0_io_a;
  wire fa_s0_c20_r0_io_b;
  wire fa_s0_c20_r0_io_ci;
  wire fa_s0_c20_r0_io_s;
  wire fa_s0_c20_r0_io_co;
  FullAdder fa_s0_c20_r0(
    .io_a(fa_s0_c20_r0_io_a),
    .io_b(fa_s0_c20_r0_io_b),
    .io_ci(fa_s0_c20_r0_io_ci),
    .io_s(fa_s0_c20_r0_io_s),
    .io_co(fa_s0_c20_r0_io_co)
  );
  wire fa_s0_c20_r1_io_a;
  wire fa_s0_c20_r1_io_b;
  wire fa_s0_c20_r1_io_ci;
  wire fa_s0_c20_r1_io_s;
  wire fa_s0_c20_r1_io_co;
  FullAdder fa_s0_c20_r1(
    .io_a(fa_s0_c20_r1_io_a),
    .io_b(fa_s0_c20_r1_io_b),
    .io_ci(fa_s0_c20_r1_io_ci),
    .io_s(fa_s0_c20_r1_io_s),
    .io_co(fa_s0_c20_r1_io_co)
  );
  wire fa_s0_c20_r2_io_a;
  wire fa_s0_c20_r2_io_b;
  wire fa_s0_c20_r2_io_ci;
  wire fa_s0_c20_r2_io_s;
  wire fa_s0_c20_r2_io_co;
  FullAdder fa_s0_c20_r2(
    .io_a(fa_s0_c20_r2_io_a),
    .io_b(fa_s0_c20_r2_io_b),
    .io_ci(fa_s0_c20_r2_io_ci),
    .io_s(fa_s0_c20_r2_io_s),
    .io_co(fa_s0_c20_r2_io_co)
  );
  wire ha_s0_c20_r3_io_a;
  wire ha_s0_c20_r3_io_b;
  wire ha_s0_c20_r3_io_s;
  wire ha_s0_c20_r3_io_co;
  HalfAdder ha_s0_c20_r3(
    .io_a(ha_s0_c20_r3_io_a),
    .io_b(ha_s0_c20_r3_io_b),
    .io_s(ha_s0_c20_r3_io_s),
    .io_co(ha_s0_c20_r3_io_co)
  );
  wire fa_s1_c20_r0_io_a;
  wire fa_s1_c20_r0_io_b;
  wire fa_s1_c20_r0_io_ci;
  wire fa_s1_c20_r0_io_s;
  wire fa_s1_c20_r0_io_co;
  FullAdder fa_s1_c20_r0(
    .io_a(fa_s1_c20_r0_io_a),
    .io_b(fa_s1_c20_r0_io_b),
    .io_ci(fa_s1_c20_r0_io_ci),
    .io_s(fa_s1_c20_r0_io_s),
    .io_co(fa_s1_c20_r0_io_co)
  );
  wire fa_s1_c20_r1_io_a;
  wire fa_s1_c20_r1_io_b;
  wire fa_s1_c20_r1_io_ci;
  wire fa_s1_c20_r1_io_s;
  wire fa_s1_c20_r1_io_co;
  FullAdder fa_s1_c20_r1(
    .io_a(fa_s1_c20_r1_io_a),
    .io_b(fa_s1_c20_r1_io_b),
    .io_ci(fa_s1_c20_r1_io_ci),
    .io_s(fa_s1_c20_r1_io_s),
    .io_co(fa_s1_c20_r1_io_co)
  );
  wire ft_s1_c20_r2_io_a;
  wire ft_s1_c20_r2_io_s;
  FallThrough ft_s1_c20_r2(
    .io_a(ft_s1_c20_r2_io_a),
    .io_s(ft_s1_c20_r2_io_s)
  );
  wire ft_s1_c20_r3_io_a;
  wire ft_s1_c20_r3_io_s;
  FallThrough ft_s1_c20_r3(
    .io_a(ft_s1_c20_r3_io_a),
    .io_s(ft_s1_c20_r3_io_s)
  );
  wire fa_s2_c20_r0_io_a;
  wire fa_s2_c20_r0_io_b;
  wire fa_s2_c20_r0_io_ci;
  wire fa_s2_c20_r0_io_s;
  wire fa_s2_c20_r0_io_co;
  FullAdder fa_s2_c20_r0(
    .io_a(fa_s2_c20_r0_io_a),
    .io_b(fa_s2_c20_r0_io_b),
    .io_ci(fa_s2_c20_r0_io_ci),
    .io_s(fa_s2_c20_r0_io_s),
    .io_co(fa_s2_c20_r0_io_co)
  );
  wire fa_s2_c20_r1_io_a;
  wire fa_s2_c20_r1_io_b;
  wire fa_s2_c20_r1_io_ci;
  wire fa_s2_c20_r1_io_s;
  wire fa_s2_c20_r1_io_co;
  FullAdder fa_s2_c20_r1(
    .io_a(fa_s2_c20_r1_io_a),
    .io_b(fa_s2_c20_r1_io_b),
    .io_ci(fa_s2_c20_r1_io_ci),
    .io_s(fa_s2_c20_r1_io_s),
    .io_co(fa_s2_c20_r1_io_co)
  );
  wire ft_s2_c20_r2_io_a;
  wire ft_s2_c20_r2_io_s;
  FallThrough ft_s2_c20_r2(
    .io_a(ft_s2_c20_r2_io_a),
    .io_s(ft_s2_c20_r2_io_s)
  );
  wire fa_s3_c20_r0_io_a;
  wire fa_s3_c20_r0_io_b;
  wire fa_s3_c20_r0_io_ci;
  wire fa_s3_c20_r0_io_s;
  wire fa_s3_c20_r0_io_co;
  FullAdder fa_s3_c20_r0(
    .io_a(fa_s3_c20_r0_io_a),
    .io_b(fa_s3_c20_r0_io_b),
    .io_ci(fa_s3_c20_r0_io_ci),
    .io_s(fa_s3_c20_r0_io_s),
    .io_co(fa_s3_c20_r0_io_co)
  );
  wire ft_s3_c20_r1_io_a;
  wire ft_s3_c20_r1_io_s;
  FallThrough ft_s3_c20_r1(
    .io_a(ft_s3_c20_r1_io_a),
    .io_s(ft_s3_c20_r1_io_s)
  );
  wire ft_s3_c20_r2_io_a;
  wire ft_s3_c20_r2_io_s;
  FallThrough ft_s3_c20_r2(
    .io_a(ft_s3_c20_r2_io_a),
    .io_s(ft_s3_c20_r2_io_s)
  );
  wire fa_s4_c20_r0_io_a;
  wire fa_s4_c20_r0_io_b;
  wire fa_s4_c20_r0_io_ci;
  wire fa_s4_c20_r0_io_s;
  wire fa_s4_c20_r0_io_co;
  FullAdder fa_s4_c20_r0(
    .io_a(fa_s4_c20_r0_io_a),
    .io_b(fa_s4_c20_r0_io_b),
    .io_ci(fa_s4_c20_r0_io_ci),
    .io_s(fa_s4_c20_r0_io_s),
    .io_co(fa_s4_c20_r0_io_co)
  );
  wire ft_s4_c20_r1_io_a;
  wire ft_s4_c20_r1_io_s;
  FallThrough ft_s4_c20_r1(
    .io_a(ft_s4_c20_r1_io_a),
    .io_s(ft_s4_c20_r1_io_s)
  );
  wire fa_s5_c20_r0_io_a;
  wire fa_s5_c20_r0_io_b;
  wire fa_s5_c20_r0_io_ci;
  wire fa_s5_c20_r0_io_s;
  wire fa_s5_c20_r0_io_co;
  FullAdder fa_s5_c20_r0(
    .io_a(fa_s5_c20_r0_io_a),
    .io_b(fa_s5_c20_r0_io_b),
    .io_ci(fa_s5_c20_r0_io_ci),
    .io_s(fa_s5_c20_r0_io_s),
    .io_co(fa_s5_c20_r0_io_co)
  );
  wire ft_s6_c20_r0_io_a;
  wire ft_s6_c20_r0_io_s;
  FallThrough ft_s6_c20_r0(
    .io_a(ft_s6_c20_r0_io_a),
    .io_s(ft_s6_c20_r0_io_s)
  );
  wire ft_s7_c20_r0_io_a;
  wire ft_s7_c20_r0_io_s;
  FallThrough ft_s7_c20_r0(
    .io_a(ft_s7_c20_r0_io_a),
    .io_s(ft_s7_c20_r0_io_s)
  );
  wire ft_s7_c20_r1_io_a;
  wire ft_s7_c20_r1_io_s;
  FallThrough ft_s7_c20_r1(
    .io_a(ft_s7_c20_r1_io_a),
    .io_s(ft_s7_c20_r1_io_s)
  );
  wire ft_s8_c20_r0_io_a;
  wire ft_s8_c20_r0_io_s;
  FallThrough ft_s8_c20_r0(
    .io_a(ft_s8_c20_r0_io_a),
    .io_s(ft_s8_c20_r0_io_s)
  );
  wire ft_s8_c20_r1_io_a;
  wire ft_s8_c20_r1_io_s;
  FallThrough ft_s8_c20_r1(
    .io_a(ft_s8_c20_r1_io_a),
    .io_s(ft_s8_c20_r1_io_s)
  );
  wire fa_s0_c21_r0_io_a;
  wire fa_s0_c21_r0_io_b;
  wire fa_s0_c21_r0_io_ci;
  wire fa_s0_c21_r0_io_s;
  wire fa_s0_c21_r0_io_co;
  FullAdder fa_s0_c21_r0(
    .io_a(fa_s0_c21_r0_io_a),
    .io_b(fa_s0_c21_r0_io_b),
    .io_ci(fa_s0_c21_r0_io_ci),
    .io_s(fa_s0_c21_r0_io_s),
    .io_co(fa_s0_c21_r0_io_co)
  );
  wire fa_s0_c21_r1_io_a;
  wire fa_s0_c21_r1_io_b;
  wire fa_s0_c21_r1_io_ci;
  wire fa_s0_c21_r1_io_s;
  wire fa_s0_c21_r1_io_co;
  FullAdder fa_s0_c21_r1(
    .io_a(fa_s0_c21_r1_io_a),
    .io_b(fa_s0_c21_r1_io_b),
    .io_ci(fa_s0_c21_r1_io_ci),
    .io_s(fa_s0_c21_r1_io_s),
    .io_co(fa_s0_c21_r1_io_co)
  );
  wire fa_s0_c21_r2_io_a;
  wire fa_s0_c21_r2_io_b;
  wire fa_s0_c21_r2_io_ci;
  wire fa_s0_c21_r2_io_s;
  wire fa_s0_c21_r2_io_co;
  FullAdder fa_s0_c21_r2(
    .io_a(fa_s0_c21_r2_io_a),
    .io_b(fa_s0_c21_r2_io_b),
    .io_ci(fa_s0_c21_r2_io_ci),
    .io_s(fa_s0_c21_r2_io_s),
    .io_co(fa_s0_c21_r2_io_co)
  );
  wire ft_s0_c21_r3_io_a;
  wire ft_s0_c21_r3_io_s;
  FallThrough ft_s0_c21_r3(
    .io_a(ft_s0_c21_r3_io_a),
    .io_s(ft_s0_c21_r3_io_s)
  );
  wire fa_s1_c21_r0_io_a;
  wire fa_s1_c21_r0_io_b;
  wire fa_s1_c21_r0_io_ci;
  wire fa_s1_c21_r0_io_s;
  wire fa_s1_c21_r0_io_co;
  FullAdder fa_s1_c21_r0(
    .io_a(fa_s1_c21_r0_io_a),
    .io_b(fa_s1_c21_r0_io_b),
    .io_ci(fa_s1_c21_r0_io_ci),
    .io_s(fa_s1_c21_r0_io_s),
    .io_co(fa_s1_c21_r0_io_co)
  );
  wire fa_s1_c21_r1_io_a;
  wire fa_s1_c21_r1_io_b;
  wire fa_s1_c21_r1_io_ci;
  wire fa_s1_c21_r1_io_s;
  wire fa_s1_c21_r1_io_co;
  FullAdder fa_s1_c21_r1(
    .io_a(fa_s1_c21_r1_io_a),
    .io_b(fa_s1_c21_r1_io_b),
    .io_ci(fa_s1_c21_r1_io_ci),
    .io_s(fa_s1_c21_r1_io_s),
    .io_co(fa_s1_c21_r1_io_co)
  );
  wire ha_s1_c21_r2_io_a;
  wire ha_s1_c21_r2_io_b;
  wire ha_s1_c21_r2_io_s;
  wire ha_s1_c21_r2_io_co;
  HalfAdder ha_s1_c21_r2(
    .io_a(ha_s1_c21_r2_io_a),
    .io_b(ha_s1_c21_r2_io_b),
    .io_s(ha_s1_c21_r2_io_s),
    .io_co(ha_s1_c21_r2_io_co)
  );
  wire fa_s2_c21_r0_io_a;
  wire fa_s2_c21_r0_io_b;
  wire fa_s2_c21_r0_io_ci;
  wire fa_s2_c21_r0_io_s;
  wire fa_s2_c21_r0_io_co;
  FullAdder fa_s2_c21_r0(
    .io_a(fa_s2_c21_r0_io_a),
    .io_b(fa_s2_c21_r0_io_b),
    .io_ci(fa_s2_c21_r0_io_ci),
    .io_s(fa_s2_c21_r0_io_s),
    .io_co(fa_s2_c21_r0_io_co)
  );
  wire ft_s2_c21_r1_io_a;
  wire ft_s2_c21_r1_io_s;
  FallThrough ft_s2_c21_r1(
    .io_a(ft_s2_c21_r1_io_a),
    .io_s(ft_s2_c21_r1_io_s)
  );
  wire ft_s2_c21_r2_io_a;
  wire ft_s2_c21_r2_io_s;
  FallThrough ft_s2_c21_r2(
    .io_a(ft_s2_c21_r2_io_a),
    .io_s(ft_s2_c21_r2_io_s)
  );
  wire fa_s3_c21_r0_io_a;
  wire fa_s3_c21_r0_io_b;
  wire fa_s3_c21_r0_io_ci;
  wire fa_s3_c21_r0_io_s;
  wire fa_s3_c21_r0_io_co;
  FullAdder fa_s3_c21_r0(
    .io_a(fa_s3_c21_r0_io_a),
    .io_b(fa_s3_c21_r0_io_b),
    .io_ci(fa_s3_c21_r0_io_ci),
    .io_s(fa_s3_c21_r0_io_s),
    .io_co(fa_s3_c21_r0_io_co)
  );
  wire ft_s3_c21_r1_io_a;
  wire ft_s3_c21_r1_io_s;
  FallThrough ft_s3_c21_r1(
    .io_a(ft_s3_c21_r1_io_a),
    .io_s(ft_s3_c21_r1_io_s)
  );
  wire ft_s3_c21_r2_io_a;
  wire ft_s3_c21_r2_io_s;
  FallThrough ft_s3_c21_r2(
    .io_a(ft_s3_c21_r2_io_a),
    .io_s(ft_s3_c21_r2_io_s)
  );
  wire fa_s4_c21_r0_io_a;
  wire fa_s4_c21_r0_io_b;
  wire fa_s4_c21_r0_io_ci;
  wire fa_s4_c21_r0_io_s;
  wire fa_s4_c21_r0_io_co;
  FullAdder fa_s4_c21_r0(
    .io_a(fa_s4_c21_r0_io_a),
    .io_b(fa_s4_c21_r0_io_b),
    .io_ci(fa_s4_c21_r0_io_ci),
    .io_s(fa_s4_c21_r0_io_s),
    .io_co(fa_s4_c21_r0_io_co)
  );
  wire ft_s4_c21_r1_io_a;
  wire ft_s4_c21_r1_io_s;
  FallThrough ft_s4_c21_r1(
    .io_a(ft_s4_c21_r1_io_a),
    .io_s(ft_s4_c21_r1_io_s)
  );
  wire fa_s5_c21_r0_io_a;
  wire fa_s5_c21_r0_io_b;
  wire fa_s5_c21_r0_io_ci;
  wire fa_s5_c21_r0_io_s;
  wire fa_s5_c21_r0_io_co;
  FullAdder fa_s5_c21_r0(
    .io_a(fa_s5_c21_r0_io_a),
    .io_b(fa_s5_c21_r0_io_b),
    .io_ci(fa_s5_c21_r0_io_ci),
    .io_s(fa_s5_c21_r0_io_s),
    .io_co(fa_s5_c21_r0_io_co)
  );
  wire ft_s6_c21_r0_io_a;
  wire ft_s6_c21_r0_io_s;
  FallThrough ft_s6_c21_r0(
    .io_a(ft_s6_c21_r0_io_a),
    .io_s(ft_s6_c21_r0_io_s)
  );
  wire ft_s6_c21_r1_io_a;
  wire ft_s6_c21_r1_io_s;
  FallThrough ft_s6_c21_r1(
    .io_a(ft_s6_c21_r1_io_a),
    .io_s(ft_s6_c21_r1_io_s)
  );
  wire ft_s7_c21_r0_io_a;
  wire ft_s7_c21_r0_io_s;
  FallThrough ft_s7_c21_r0(
    .io_a(ft_s7_c21_r0_io_a),
    .io_s(ft_s7_c21_r0_io_s)
  );
  wire ft_s7_c21_r1_io_a;
  wire ft_s7_c21_r1_io_s;
  FallThrough ft_s7_c21_r1(
    .io_a(ft_s7_c21_r1_io_a),
    .io_s(ft_s7_c21_r1_io_s)
  );
  wire ft_s8_c21_r0_io_a;
  wire ft_s8_c21_r0_io_s;
  FallThrough ft_s8_c21_r0(
    .io_a(ft_s8_c21_r0_io_a),
    .io_s(ft_s8_c21_r0_io_s)
  );
  wire ft_s8_c21_r1_io_a;
  wire ft_s8_c21_r1_io_s;
  FallThrough ft_s8_c21_r1(
    .io_a(ft_s8_c21_r1_io_a),
    .io_s(ft_s8_c21_r1_io_s)
  );
  wire fa_s0_c22_r0_io_a;
  wire fa_s0_c22_r0_io_b;
  wire fa_s0_c22_r0_io_ci;
  wire fa_s0_c22_r0_io_s;
  wire fa_s0_c22_r0_io_co;
  FullAdder fa_s0_c22_r0(
    .io_a(fa_s0_c22_r0_io_a),
    .io_b(fa_s0_c22_r0_io_b),
    .io_ci(fa_s0_c22_r0_io_ci),
    .io_s(fa_s0_c22_r0_io_s),
    .io_co(fa_s0_c22_r0_io_co)
  );
  wire fa_s0_c22_r1_io_a;
  wire fa_s0_c22_r1_io_b;
  wire fa_s0_c22_r1_io_ci;
  wire fa_s0_c22_r1_io_s;
  wire fa_s0_c22_r1_io_co;
  FullAdder fa_s0_c22_r1(
    .io_a(fa_s0_c22_r1_io_a),
    .io_b(fa_s0_c22_r1_io_b),
    .io_ci(fa_s0_c22_r1_io_ci),
    .io_s(fa_s0_c22_r1_io_s),
    .io_co(fa_s0_c22_r1_io_co)
  );
  wire fa_s0_c22_r2_io_a;
  wire fa_s0_c22_r2_io_b;
  wire fa_s0_c22_r2_io_ci;
  wire fa_s0_c22_r2_io_s;
  wire fa_s0_c22_r2_io_co;
  FullAdder fa_s0_c22_r2(
    .io_a(fa_s0_c22_r2_io_a),
    .io_b(fa_s0_c22_r2_io_b),
    .io_ci(fa_s0_c22_r2_io_ci),
    .io_s(fa_s0_c22_r2_io_s),
    .io_co(fa_s0_c22_r2_io_co)
  );
  wire fa_s1_c22_r0_io_a;
  wire fa_s1_c22_r0_io_b;
  wire fa_s1_c22_r0_io_ci;
  wire fa_s1_c22_r0_io_s;
  wire fa_s1_c22_r0_io_co;
  FullAdder fa_s1_c22_r0(
    .io_a(fa_s1_c22_r0_io_a),
    .io_b(fa_s1_c22_r0_io_b),
    .io_ci(fa_s1_c22_r0_io_ci),
    .io_s(fa_s1_c22_r0_io_s),
    .io_co(fa_s1_c22_r0_io_co)
  );
  wire fa_s1_c22_r1_io_a;
  wire fa_s1_c22_r1_io_b;
  wire fa_s1_c22_r1_io_ci;
  wire fa_s1_c22_r1_io_s;
  wire fa_s1_c22_r1_io_co;
  FullAdder fa_s1_c22_r1(
    .io_a(fa_s1_c22_r1_io_a),
    .io_b(fa_s1_c22_r1_io_b),
    .io_ci(fa_s1_c22_r1_io_ci),
    .io_s(fa_s1_c22_r1_io_s),
    .io_co(fa_s1_c22_r1_io_co)
  );
  wire fa_s2_c22_r0_io_a;
  wire fa_s2_c22_r0_io_b;
  wire fa_s2_c22_r0_io_ci;
  wire fa_s2_c22_r0_io_s;
  wire fa_s2_c22_r0_io_co;
  FullAdder fa_s2_c22_r0(
    .io_a(fa_s2_c22_r0_io_a),
    .io_b(fa_s2_c22_r0_io_b),
    .io_ci(fa_s2_c22_r0_io_ci),
    .io_s(fa_s2_c22_r0_io_s),
    .io_co(fa_s2_c22_r0_io_co)
  );
  wire ha_s2_c22_r1_io_a;
  wire ha_s2_c22_r1_io_b;
  wire ha_s2_c22_r1_io_s;
  wire ha_s2_c22_r1_io_co;
  HalfAdder ha_s2_c22_r1(
    .io_a(ha_s2_c22_r1_io_a),
    .io_b(ha_s2_c22_r1_io_b),
    .io_s(ha_s2_c22_r1_io_s),
    .io_co(ha_s2_c22_r1_io_co)
  );
  wire fa_s3_c22_r0_io_a;
  wire fa_s3_c22_r0_io_b;
  wire fa_s3_c22_r0_io_ci;
  wire fa_s3_c22_r0_io_s;
  wire fa_s3_c22_r0_io_co;
  FullAdder fa_s3_c22_r0(
    .io_a(fa_s3_c22_r0_io_a),
    .io_b(fa_s3_c22_r0_io_b),
    .io_ci(fa_s3_c22_r0_io_ci),
    .io_s(fa_s3_c22_r0_io_s),
    .io_co(fa_s3_c22_r0_io_co)
  );
  wire ft_s4_c22_r0_io_a;
  wire ft_s4_c22_r0_io_s;
  FallThrough ft_s4_c22_r0(
    .io_a(ft_s4_c22_r0_io_a),
    .io_s(ft_s4_c22_r0_io_s)
  );
  wire ft_s4_c22_r1_io_a;
  wire ft_s4_c22_r1_io_s;
  FallThrough ft_s4_c22_r1(
    .io_a(ft_s4_c22_r1_io_a),
    .io_s(ft_s4_c22_r1_io_s)
  );
  wire fa_s5_c22_r0_io_a;
  wire fa_s5_c22_r0_io_b;
  wire fa_s5_c22_r0_io_ci;
  wire fa_s5_c22_r0_io_s;
  wire fa_s5_c22_r0_io_co;
  FullAdder fa_s5_c22_r0(
    .io_a(fa_s5_c22_r0_io_a),
    .io_b(fa_s5_c22_r0_io_b),
    .io_ci(fa_s5_c22_r0_io_ci),
    .io_s(fa_s5_c22_r0_io_s),
    .io_co(fa_s5_c22_r0_io_co)
  );
  wire ft_s6_c22_r0_io_a;
  wire ft_s6_c22_r0_io_s;
  FallThrough ft_s6_c22_r0(
    .io_a(ft_s6_c22_r0_io_a),
    .io_s(ft_s6_c22_r0_io_s)
  );
  wire ft_s6_c22_r1_io_a;
  wire ft_s6_c22_r1_io_s;
  FallThrough ft_s6_c22_r1(
    .io_a(ft_s6_c22_r1_io_a),
    .io_s(ft_s6_c22_r1_io_s)
  );
  wire ft_s7_c22_r0_io_a;
  wire ft_s7_c22_r0_io_s;
  FallThrough ft_s7_c22_r0(
    .io_a(ft_s7_c22_r0_io_a),
    .io_s(ft_s7_c22_r0_io_s)
  );
  wire ft_s7_c22_r1_io_a;
  wire ft_s7_c22_r1_io_s;
  FallThrough ft_s7_c22_r1(
    .io_a(ft_s7_c22_r1_io_a),
    .io_s(ft_s7_c22_r1_io_s)
  );
  wire ft_s8_c22_r0_io_a;
  wire ft_s8_c22_r0_io_s;
  FallThrough ft_s8_c22_r0(
    .io_a(ft_s8_c22_r0_io_a),
    .io_s(ft_s8_c22_r0_io_s)
  );
  wire ft_s8_c22_r1_io_a;
  wire ft_s8_c22_r1_io_s;
  FallThrough ft_s8_c22_r1(
    .io_a(ft_s8_c22_r1_io_a),
    .io_s(ft_s8_c22_r1_io_s)
  );
  wire fa_s0_c23_r0_io_a;
  wire fa_s0_c23_r0_io_b;
  wire fa_s0_c23_r0_io_ci;
  wire fa_s0_c23_r0_io_s;
  wire fa_s0_c23_r0_io_co;
  FullAdder fa_s0_c23_r0(
    .io_a(fa_s0_c23_r0_io_a),
    .io_b(fa_s0_c23_r0_io_b),
    .io_ci(fa_s0_c23_r0_io_ci),
    .io_s(fa_s0_c23_r0_io_s),
    .io_co(fa_s0_c23_r0_io_co)
  );
  wire fa_s0_c23_r1_io_a;
  wire fa_s0_c23_r1_io_b;
  wire fa_s0_c23_r1_io_ci;
  wire fa_s0_c23_r1_io_s;
  wire fa_s0_c23_r1_io_co;
  FullAdder fa_s0_c23_r1(
    .io_a(fa_s0_c23_r1_io_a),
    .io_b(fa_s0_c23_r1_io_b),
    .io_ci(fa_s0_c23_r1_io_ci),
    .io_s(fa_s0_c23_r1_io_s),
    .io_co(fa_s0_c23_r1_io_co)
  );
  wire ft_s0_c23_r2_io_a;
  wire ft_s0_c23_r2_io_s;
  FallThrough ft_s0_c23_r2(
    .io_a(ft_s0_c23_r2_io_a),
    .io_s(ft_s0_c23_r2_io_s)
  );
  wire ft_s0_c23_r3_io_a;
  wire ft_s0_c23_r3_io_s;
  FallThrough ft_s0_c23_r3(
    .io_a(ft_s0_c23_r3_io_a),
    .io_s(ft_s0_c23_r3_io_s)
  );
  wire fa_s1_c23_r0_io_a;
  wire fa_s1_c23_r0_io_b;
  wire fa_s1_c23_r0_io_ci;
  wire fa_s1_c23_r0_io_s;
  wire fa_s1_c23_r0_io_co;
  FullAdder fa_s1_c23_r0(
    .io_a(fa_s1_c23_r0_io_a),
    .io_b(fa_s1_c23_r0_io_b),
    .io_ci(fa_s1_c23_r0_io_ci),
    .io_s(fa_s1_c23_r0_io_s),
    .io_co(fa_s1_c23_r0_io_co)
  );
  wire fa_s1_c23_r1_io_a;
  wire fa_s1_c23_r1_io_b;
  wire fa_s1_c23_r1_io_ci;
  wire fa_s1_c23_r1_io_s;
  wire fa_s1_c23_r1_io_co;
  FullAdder fa_s1_c23_r1(
    .io_a(fa_s1_c23_r1_io_a),
    .io_b(fa_s1_c23_r1_io_b),
    .io_ci(fa_s1_c23_r1_io_ci),
    .io_s(fa_s1_c23_r1_io_s),
    .io_co(fa_s1_c23_r1_io_co)
  );
  wire ft_s1_c23_r2_io_a;
  wire ft_s1_c23_r2_io_s;
  FallThrough ft_s1_c23_r2(
    .io_a(ft_s1_c23_r2_io_a),
    .io_s(ft_s1_c23_r2_io_s)
  );
  wire fa_s2_c23_r0_io_a;
  wire fa_s2_c23_r0_io_b;
  wire fa_s2_c23_r0_io_ci;
  wire fa_s2_c23_r0_io_s;
  wire fa_s2_c23_r0_io_co;
  FullAdder fa_s2_c23_r0(
    .io_a(fa_s2_c23_r0_io_a),
    .io_b(fa_s2_c23_r0_io_b),
    .io_ci(fa_s2_c23_r0_io_ci),
    .io_s(fa_s2_c23_r0_io_s),
    .io_co(fa_s2_c23_r0_io_co)
  );
  wire ft_s2_c23_r1_io_a;
  wire ft_s2_c23_r1_io_s;
  FallThrough ft_s2_c23_r1(
    .io_a(ft_s2_c23_r1_io_a),
    .io_s(ft_s2_c23_r1_io_s)
  );
  wire ft_s2_c23_r2_io_a;
  wire ft_s2_c23_r2_io_s;
  FallThrough ft_s2_c23_r2(
    .io_a(ft_s2_c23_r2_io_a),
    .io_s(ft_s2_c23_r2_io_s)
  );
  wire fa_s3_c23_r0_io_a;
  wire fa_s3_c23_r0_io_b;
  wire fa_s3_c23_r0_io_ci;
  wire fa_s3_c23_r0_io_s;
  wire fa_s3_c23_r0_io_co;
  FullAdder fa_s3_c23_r0(
    .io_a(fa_s3_c23_r0_io_a),
    .io_b(fa_s3_c23_r0_io_b),
    .io_ci(fa_s3_c23_r0_io_ci),
    .io_s(fa_s3_c23_r0_io_s),
    .io_co(fa_s3_c23_r0_io_co)
  );
  wire ft_s3_c23_r1_io_a;
  wire ft_s3_c23_r1_io_s;
  FallThrough ft_s3_c23_r1(
    .io_a(ft_s3_c23_r1_io_a),
    .io_s(ft_s3_c23_r1_io_s)
  );
  wire ft_s3_c23_r2_io_a;
  wire ft_s3_c23_r2_io_s;
  FallThrough ft_s3_c23_r2(
    .io_a(ft_s3_c23_r2_io_a),
    .io_s(ft_s3_c23_r2_io_s)
  );
  wire fa_s4_c23_r0_io_a;
  wire fa_s4_c23_r0_io_b;
  wire fa_s4_c23_r0_io_ci;
  wire fa_s4_c23_r0_io_s;
  wire fa_s4_c23_r0_io_co;
  FullAdder fa_s4_c23_r0(
    .io_a(fa_s4_c23_r0_io_a),
    .io_b(fa_s4_c23_r0_io_b),
    .io_ci(fa_s4_c23_r0_io_ci),
    .io_s(fa_s4_c23_r0_io_s),
    .io_co(fa_s4_c23_r0_io_co)
  );
  wire ft_s4_c23_r1_io_a;
  wire ft_s4_c23_r1_io_s;
  FallThrough ft_s4_c23_r1(
    .io_a(ft_s4_c23_r1_io_a),
    .io_s(ft_s4_c23_r1_io_s)
  );
  wire ft_s5_c23_r0_io_a;
  wire ft_s5_c23_r0_io_s;
  FallThrough ft_s5_c23_r0(
    .io_a(ft_s5_c23_r0_io_a),
    .io_s(ft_s5_c23_r0_io_s)
  );
  wire ft_s5_c23_r1_io_a;
  wire ft_s5_c23_r1_io_s;
  FallThrough ft_s5_c23_r1(
    .io_a(ft_s5_c23_r1_io_a),
    .io_s(ft_s5_c23_r1_io_s)
  );
  wire fa_s6_c23_r0_io_a;
  wire fa_s6_c23_r0_io_b;
  wire fa_s6_c23_r0_io_ci;
  wire fa_s6_c23_r0_io_s;
  wire fa_s6_c23_r0_io_co;
  FullAdder fa_s6_c23_r0(
    .io_a(fa_s6_c23_r0_io_a),
    .io_b(fa_s6_c23_r0_io_b),
    .io_ci(fa_s6_c23_r0_io_ci),
    .io_s(fa_s6_c23_r0_io_s),
    .io_co(fa_s6_c23_r0_io_co)
  );
  wire ft_s7_c23_r0_io_a;
  wire ft_s7_c23_r0_io_s;
  FallThrough ft_s7_c23_r0(
    .io_a(ft_s7_c23_r0_io_a),
    .io_s(ft_s7_c23_r0_io_s)
  );
  wire ft_s8_c23_r0_io_a;
  wire ft_s8_c23_r0_io_s;
  FallThrough ft_s8_c23_r0(
    .io_a(ft_s8_c23_r0_io_a),
    .io_s(ft_s8_c23_r0_io_s)
  );
  wire fa_s0_c24_r0_io_a;
  wire fa_s0_c24_r0_io_b;
  wire fa_s0_c24_r0_io_ci;
  wire fa_s0_c24_r0_io_s;
  wire fa_s0_c24_r0_io_co;
  FullAdder fa_s0_c24_r0(
    .io_a(fa_s0_c24_r0_io_a),
    .io_b(fa_s0_c24_r0_io_b),
    .io_ci(fa_s0_c24_r0_io_ci),
    .io_s(fa_s0_c24_r0_io_s),
    .io_co(fa_s0_c24_r0_io_co)
  );
  wire fa_s0_c24_r1_io_a;
  wire fa_s0_c24_r1_io_b;
  wire fa_s0_c24_r1_io_ci;
  wire fa_s0_c24_r1_io_s;
  wire fa_s0_c24_r1_io_co;
  FullAdder fa_s0_c24_r1(
    .io_a(fa_s0_c24_r1_io_a),
    .io_b(fa_s0_c24_r1_io_b),
    .io_ci(fa_s0_c24_r1_io_ci),
    .io_s(fa_s0_c24_r1_io_s),
    .io_co(fa_s0_c24_r1_io_co)
  );
  wire ft_s0_c24_r2_io_a;
  wire ft_s0_c24_r2_io_s;
  FallThrough ft_s0_c24_r2(
    .io_a(ft_s0_c24_r2_io_a),
    .io_s(ft_s0_c24_r2_io_s)
  );
  wire fa_s1_c24_r0_io_a;
  wire fa_s1_c24_r0_io_b;
  wire fa_s1_c24_r0_io_ci;
  wire fa_s1_c24_r0_io_s;
  wire fa_s1_c24_r0_io_co;
  FullAdder fa_s1_c24_r0(
    .io_a(fa_s1_c24_r0_io_a),
    .io_b(fa_s1_c24_r0_io_b),
    .io_ci(fa_s1_c24_r0_io_ci),
    .io_s(fa_s1_c24_r0_io_s),
    .io_co(fa_s1_c24_r0_io_co)
  );
  wire ft_s1_c24_r1_io_a;
  wire ft_s1_c24_r1_io_s;
  FallThrough ft_s1_c24_r1(
    .io_a(ft_s1_c24_r1_io_a),
    .io_s(ft_s1_c24_r1_io_s)
  );
  wire ft_s1_c24_r2_io_a;
  wire ft_s1_c24_r2_io_s;
  FallThrough ft_s1_c24_r2(
    .io_a(ft_s1_c24_r2_io_a),
    .io_s(ft_s1_c24_r2_io_s)
  );
  wire fa_s2_c24_r0_io_a;
  wire fa_s2_c24_r0_io_b;
  wire fa_s2_c24_r0_io_ci;
  wire fa_s2_c24_r0_io_s;
  wire fa_s2_c24_r0_io_co;
  FullAdder fa_s2_c24_r0(
    .io_a(fa_s2_c24_r0_io_a),
    .io_b(fa_s2_c24_r0_io_b),
    .io_ci(fa_s2_c24_r0_io_ci),
    .io_s(fa_s2_c24_r0_io_s),
    .io_co(fa_s2_c24_r0_io_co)
  );
  wire ft_s2_c24_r1_io_a;
  wire ft_s2_c24_r1_io_s;
  FallThrough ft_s2_c24_r1(
    .io_a(ft_s2_c24_r1_io_a),
    .io_s(ft_s2_c24_r1_io_s)
  );
  wire ft_s2_c24_r2_io_a;
  wire ft_s2_c24_r2_io_s;
  FallThrough ft_s2_c24_r2(
    .io_a(ft_s2_c24_r2_io_a),
    .io_s(ft_s2_c24_r2_io_s)
  );
  wire fa_s3_c24_r0_io_a;
  wire fa_s3_c24_r0_io_b;
  wire fa_s3_c24_r0_io_ci;
  wire fa_s3_c24_r0_io_s;
  wire fa_s3_c24_r0_io_co;
  FullAdder fa_s3_c24_r0(
    .io_a(fa_s3_c24_r0_io_a),
    .io_b(fa_s3_c24_r0_io_b),
    .io_ci(fa_s3_c24_r0_io_ci),
    .io_s(fa_s3_c24_r0_io_s),
    .io_co(fa_s3_c24_r0_io_co)
  );
  wire ft_s3_c24_r1_io_a;
  wire ft_s3_c24_r1_io_s;
  FallThrough ft_s3_c24_r1(
    .io_a(ft_s3_c24_r1_io_a),
    .io_s(ft_s3_c24_r1_io_s)
  );
  wire fa_s4_c24_r0_io_a;
  wire fa_s4_c24_r0_io_b;
  wire fa_s4_c24_r0_io_ci;
  wire fa_s4_c24_r0_io_s;
  wire fa_s4_c24_r0_io_co;
  FullAdder fa_s4_c24_r0(
    .io_a(fa_s4_c24_r0_io_a),
    .io_b(fa_s4_c24_r0_io_b),
    .io_ci(fa_s4_c24_r0_io_ci),
    .io_s(fa_s4_c24_r0_io_s),
    .io_co(fa_s4_c24_r0_io_co)
  );
  wire ft_s5_c24_r0_io_a;
  wire ft_s5_c24_r0_io_s;
  FallThrough ft_s5_c24_r0(
    .io_a(ft_s5_c24_r0_io_a),
    .io_s(ft_s5_c24_r0_io_s)
  );
  wire ft_s5_c24_r1_io_a;
  wire ft_s5_c24_r1_io_s;
  FallThrough ft_s5_c24_r1(
    .io_a(ft_s5_c24_r1_io_a),
    .io_s(ft_s5_c24_r1_io_s)
  );
  wire ft_s6_c24_r0_io_a;
  wire ft_s6_c24_r0_io_s;
  FallThrough ft_s6_c24_r0(
    .io_a(ft_s6_c24_r0_io_a),
    .io_s(ft_s6_c24_r0_io_s)
  );
  wire ft_s6_c24_r1_io_a;
  wire ft_s6_c24_r1_io_s;
  FallThrough ft_s6_c24_r1(
    .io_a(ft_s6_c24_r1_io_a),
    .io_s(ft_s6_c24_r1_io_s)
  );
  wire fa_s7_c24_r0_io_a;
  wire fa_s7_c24_r0_io_b;
  wire fa_s7_c24_r0_io_ci;
  wire fa_s7_c24_r0_io_s;
  wire fa_s7_c24_r0_io_co;
  FullAdder fa_s7_c24_r0(
    .io_a(fa_s7_c24_r0_io_a),
    .io_b(fa_s7_c24_r0_io_b),
    .io_ci(fa_s7_c24_r0_io_ci),
    .io_s(fa_s7_c24_r0_io_s),
    .io_co(fa_s7_c24_r0_io_co)
  );
  wire ft_s8_c24_r0_io_a;
  wire ft_s8_c24_r0_io_s;
  FallThrough ft_s8_c24_r0(
    .io_a(ft_s8_c24_r0_io_a),
    .io_s(ft_s8_c24_r0_io_s)
  );
  wire fa_s0_c25_r0_io_a;
  wire fa_s0_c25_r0_io_b;
  wire fa_s0_c25_r0_io_ci;
  wire fa_s0_c25_r0_io_s;
  wire fa_s0_c25_r0_io_co;
  FullAdder fa_s0_c25_r0(
    .io_a(fa_s0_c25_r0_io_a),
    .io_b(fa_s0_c25_r0_io_b),
    .io_ci(fa_s0_c25_r0_io_ci),
    .io_s(fa_s0_c25_r0_io_s),
    .io_co(fa_s0_c25_r0_io_co)
  );
  wire fa_s0_c25_r1_io_a;
  wire fa_s0_c25_r1_io_b;
  wire fa_s0_c25_r1_io_ci;
  wire fa_s0_c25_r1_io_s;
  wire fa_s0_c25_r1_io_co;
  FullAdder fa_s0_c25_r1(
    .io_a(fa_s0_c25_r1_io_a),
    .io_b(fa_s0_c25_r1_io_b),
    .io_ci(fa_s0_c25_r1_io_ci),
    .io_s(fa_s0_c25_r1_io_s),
    .io_co(fa_s0_c25_r1_io_co)
  );
  wire fa_s1_c25_r0_io_a;
  wire fa_s1_c25_r0_io_b;
  wire fa_s1_c25_r0_io_ci;
  wire fa_s1_c25_r0_io_s;
  wire fa_s1_c25_r0_io_co;
  FullAdder fa_s1_c25_r0(
    .io_a(fa_s1_c25_r0_io_a),
    .io_b(fa_s1_c25_r0_io_b),
    .io_ci(fa_s1_c25_r0_io_ci),
    .io_s(fa_s1_c25_r0_io_s),
    .io_co(fa_s1_c25_r0_io_co)
  );
  wire ft_s1_c25_r1_io_a;
  wire ft_s1_c25_r1_io_s;
  FallThrough ft_s1_c25_r1(
    .io_a(ft_s1_c25_r1_io_a),
    .io_s(ft_s1_c25_r1_io_s)
  );
  wire fa_s2_c25_r0_io_a;
  wire fa_s2_c25_r0_io_b;
  wire fa_s2_c25_r0_io_ci;
  wire fa_s2_c25_r0_io_s;
  wire fa_s2_c25_r0_io_co;
  FullAdder fa_s2_c25_r0(
    .io_a(fa_s2_c25_r0_io_a),
    .io_b(fa_s2_c25_r0_io_b),
    .io_ci(fa_s2_c25_r0_io_ci),
    .io_s(fa_s2_c25_r0_io_s),
    .io_co(fa_s2_c25_r0_io_co)
  );
  wire ha_s3_c25_r0_io_a;
  wire ha_s3_c25_r0_io_b;
  wire ha_s3_c25_r0_io_s;
  wire ha_s3_c25_r0_io_co;
  HalfAdder ha_s3_c25_r0(
    .io_a(ha_s3_c25_r0_io_a),
    .io_b(ha_s3_c25_r0_io_b),
    .io_s(ha_s3_c25_r0_io_s),
    .io_co(ha_s3_c25_r0_io_co)
  );
  wire ha_s4_c25_r0_io_a;
  wire ha_s4_c25_r0_io_b;
  wire ha_s4_c25_r0_io_s;
  wire ha_s4_c25_r0_io_co;
  HalfAdder ha_s4_c25_r0(
    .io_a(ha_s4_c25_r0_io_a),
    .io_b(ha_s4_c25_r0_io_b),
    .io_s(ha_s4_c25_r0_io_s),
    .io_co(ha_s4_c25_r0_io_co)
  );
  wire ft_s5_c25_r0_io_a;
  wire ft_s5_c25_r0_io_s;
  FallThrough ft_s5_c25_r0(
    .io_a(ft_s5_c25_r0_io_a),
    .io_s(ft_s5_c25_r0_io_s)
  );
  wire ft_s5_c25_r1_io_a;
  wire ft_s5_c25_r1_io_s;
  FallThrough ft_s5_c25_r1(
    .io_a(ft_s5_c25_r1_io_a),
    .io_s(ft_s5_c25_r1_io_s)
  );
  wire ft_s6_c25_r0_io_a;
  wire ft_s6_c25_r0_io_s;
  FallThrough ft_s6_c25_r0(
    .io_a(ft_s6_c25_r0_io_a),
    .io_s(ft_s6_c25_r0_io_s)
  );
  wire ft_s6_c25_r1_io_a;
  wire ft_s6_c25_r1_io_s;
  FallThrough ft_s6_c25_r1(
    .io_a(ft_s6_c25_r1_io_a),
    .io_s(ft_s6_c25_r1_io_s)
  );
  wire ft_s7_c25_r0_io_a;
  wire ft_s7_c25_r0_io_s;
  FallThrough ft_s7_c25_r0(
    .io_a(ft_s7_c25_r0_io_a),
    .io_s(ft_s7_c25_r0_io_s)
  );
  wire ft_s7_c25_r1_io_a;
  wire ft_s7_c25_r1_io_s;
  FallThrough ft_s7_c25_r1(
    .io_a(ft_s7_c25_r1_io_a),
    .io_s(ft_s7_c25_r1_io_s)
  );
  wire fa_s8_c25_r0_io_a;
  wire fa_s8_c25_r0_io_b;
  wire fa_s8_c25_r0_io_ci;
  wire fa_s8_c25_r0_io_s;
  wire fa_s8_c25_r0_io_co;
  FullAdder fa_s8_c25_r0(
    .io_a(fa_s8_c25_r0_io_a),
    .io_b(fa_s8_c25_r0_io_b),
    .io_ci(fa_s8_c25_r0_io_ci),
    .io_s(fa_s8_c25_r0_io_s),
    .io_co(fa_s8_c25_r0_io_co)
  );
  wire fa_s0_c26_r0_io_a;
  wire fa_s0_c26_r0_io_b;
  wire fa_s0_c26_r0_io_ci;
  wire fa_s0_c26_r0_io_s;
  wire fa_s0_c26_r0_io_co;
  FullAdder fa_s0_c26_r0(
    .io_a(fa_s0_c26_r0_io_a),
    .io_b(fa_s0_c26_r0_io_b),
    .io_ci(fa_s0_c26_r0_io_ci),
    .io_s(fa_s0_c26_r0_io_s),
    .io_co(fa_s0_c26_r0_io_co)
  );
  wire ft_s0_c26_r1_io_a;
  wire ft_s0_c26_r1_io_s;
  FallThrough ft_s0_c26_r1(
    .io_a(ft_s0_c26_r1_io_a),
    .io_s(ft_s0_c26_r1_io_s)
  );
  wire ft_s0_c26_r2_io_a;
  wire ft_s0_c26_r2_io_s;
  FallThrough ft_s0_c26_r2(
    .io_a(ft_s0_c26_r2_io_a),
    .io_s(ft_s0_c26_r2_io_s)
  );
  wire fa_s1_c26_r0_io_a;
  wire fa_s1_c26_r0_io_b;
  wire fa_s1_c26_r0_io_ci;
  wire fa_s1_c26_r0_io_s;
  wire fa_s1_c26_r0_io_co;
  FullAdder fa_s1_c26_r0(
    .io_a(fa_s1_c26_r0_io_a),
    .io_b(fa_s1_c26_r0_io_b),
    .io_ci(fa_s1_c26_r0_io_ci),
    .io_s(fa_s1_c26_r0_io_s),
    .io_co(fa_s1_c26_r0_io_co)
  );
  wire ft_s1_c26_r1_io_a;
  wire ft_s1_c26_r1_io_s;
  FallThrough ft_s1_c26_r1(
    .io_a(ft_s1_c26_r1_io_a),
    .io_s(ft_s1_c26_r1_io_s)
  );
  wire ft_s1_c26_r2_io_a;
  wire ft_s1_c26_r2_io_s;
  FallThrough ft_s1_c26_r2(
    .io_a(ft_s1_c26_r2_io_a),
    .io_s(ft_s1_c26_r2_io_s)
  );
  wire fa_s2_c26_r0_io_a;
  wire fa_s2_c26_r0_io_b;
  wire fa_s2_c26_r0_io_ci;
  wire fa_s2_c26_r0_io_s;
  wire fa_s2_c26_r0_io_co;
  FullAdder fa_s2_c26_r0(
    .io_a(fa_s2_c26_r0_io_a),
    .io_b(fa_s2_c26_r0_io_b),
    .io_ci(fa_s2_c26_r0_io_ci),
    .io_s(fa_s2_c26_r0_io_s),
    .io_co(fa_s2_c26_r0_io_co)
  );
  wire ft_s2_c26_r1_io_a;
  wire ft_s2_c26_r1_io_s;
  FallThrough ft_s2_c26_r1(
    .io_a(ft_s2_c26_r1_io_a),
    .io_s(ft_s2_c26_r1_io_s)
  );
  wire fa_s3_c26_r0_io_a;
  wire fa_s3_c26_r0_io_b;
  wire fa_s3_c26_r0_io_ci;
  wire fa_s3_c26_r0_io_s;
  wire fa_s3_c26_r0_io_co;
  FullAdder fa_s3_c26_r0(
    .io_a(fa_s3_c26_r0_io_a),
    .io_b(fa_s3_c26_r0_io_b),
    .io_ci(fa_s3_c26_r0_io_ci),
    .io_s(fa_s3_c26_r0_io_s),
    .io_co(fa_s3_c26_r0_io_co)
  );
  wire ft_s4_c26_r0_io_a;
  wire ft_s4_c26_r0_io_s;
  FallThrough ft_s4_c26_r0(
    .io_a(ft_s4_c26_r0_io_a),
    .io_s(ft_s4_c26_r0_io_s)
  );
  wire ft_s4_c26_r1_io_a;
  wire ft_s4_c26_r1_io_s;
  FallThrough ft_s4_c26_r1(
    .io_a(ft_s4_c26_r1_io_a),
    .io_s(ft_s4_c26_r1_io_s)
  );
  wire fa_s5_c26_r0_io_a;
  wire fa_s5_c26_r0_io_b;
  wire fa_s5_c26_r0_io_ci;
  wire fa_s5_c26_r0_io_s;
  wire fa_s5_c26_r0_io_co;
  FullAdder fa_s5_c26_r0(
    .io_a(fa_s5_c26_r0_io_a),
    .io_b(fa_s5_c26_r0_io_b),
    .io_ci(fa_s5_c26_r0_io_ci),
    .io_s(fa_s5_c26_r0_io_s),
    .io_co(fa_s5_c26_r0_io_co)
  );
  wire ft_s6_c26_r0_io_a;
  wire ft_s6_c26_r0_io_s;
  FallThrough ft_s6_c26_r0(
    .io_a(ft_s6_c26_r0_io_a),
    .io_s(ft_s6_c26_r0_io_s)
  );
  wire ft_s7_c26_r0_io_a;
  wire ft_s7_c26_r0_io_s;
  FallThrough ft_s7_c26_r0(
    .io_a(ft_s7_c26_r0_io_a),
    .io_s(ft_s7_c26_r0_io_s)
  );
  wire ft_s8_c26_r0_io_a;
  wire ft_s8_c26_r0_io_s;
  FallThrough ft_s8_c26_r0(
    .io_a(ft_s8_c26_r0_io_a),
    .io_s(ft_s8_c26_r0_io_s)
  );
  wire fa_s0_c27_r0_io_a;
  wire fa_s0_c27_r0_io_b;
  wire fa_s0_c27_r0_io_ci;
  wire fa_s0_c27_r0_io_s;
  wire fa_s0_c27_r0_io_co;
  FullAdder fa_s0_c27_r0(
    .io_a(fa_s0_c27_r0_io_a),
    .io_b(fa_s0_c27_r0_io_b),
    .io_ci(fa_s0_c27_r0_io_ci),
    .io_s(fa_s0_c27_r0_io_s),
    .io_co(fa_s0_c27_r0_io_co)
  );
  wire ft_s0_c27_r1_io_a;
  wire ft_s0_c27_r1_io_s;
  FallThrough ft_s0_c27_r1(
    .io_a(ft_s0_c27_r1_io_a),
    .io_s(ft_s0_c27_r1_io_s)
  );
  wire fa_s1_c27_r0_io_a;
  wire fa_s1_c27_r0_io_b;
  wire fa_s1_c27_r0_io_ci;
  wire fa_s1_c27_r0_io_s;
  wire fa_s1_c27_r0_io_co;
  FullAdder fa_s1_c27_r0(
    .io_a(fa_s1_c27_r0_io_a),
    .io_b(fa_s1_c27_r0_io_b),
    .io_ci(fa_s1_c27_r0_io_ci),
    .io_s(fa_s1_c27_r0_io_s),
    .io_co(fa_s1_c27_r0_io_co)
  );
  wire ft_s2_c27_r0_io_a;
  wire ft_s2_c27_r0_io_s;
  FallThrough ft_s2_c27_r0(
    .io_a(ft_s2_c27_r0_io_a),
    .io_s(ft_s2_c27_r0_io_s)
  );
  wire ft_s2_c27_r1_io_a;
  wire ft_s2_c27_r1_io_s;
  FallThrough ft_s2_c27_r1(
    .io_a(ft_s2_c27_r1_io_a),
    .io_s(ft_s2_c27_r1_io_s)
  );
  wire fa_s3_c27_r0_io_a;
  wire fa_s3_c27_r0_io_b;
  wire fa_s3_c27_r0_io_ci;
  wire fa_s3_c27_r0_io_s;
  wire fa_s3_c27_r0_io_co;
  FullAdder fa_s3_c27_r0(
    .io_a(fa_s3_c27_r0_io_a),
    .io_b(fa_s3_c27_r0_io_b),
    .io_ci(fa_s3_c27_r0_io_ci),
    .io_s(fa_s3_c27_r0_io_s),
    .io_co(fa_s3_c27_r0_io_co)
  );
  wire ft_s4_c27_r0_io_a;
  wire ft_s4_c27_r0_io_s;
  FallThrough ft_s4_c27_r0(
    .io_a(ft_s4_c27_r0_io_a),
    .io_s(ft_s4_c27_r0_io_s)
  );
  wire ft_s4_c27_r1_io_a;
  wire ft_s4_c27_r1_io_s;
  FallThrough ft_s4_c27_r1(
    .io_a(ft_s4_c27_r1_io_a),
    .io_s(ft_s4_c27_r1_io_s)
  );
  wire ft_s5_c27_r0_io_a;
  wire ft_s5_c27_r0_io_s;
  FallThrough ft_s5_c27_r0(
    .io_a(ft_s5_c27_r0_io_a),
    .io_s(ft_s5_c27_r0_io_s)
  );
  wire ft_s5_c27_r1_io_a;
  wire ft_s5_c27_r1_io_s;
  FallThrough ft_s5_c27_r1(
    .io_a(ft_s5_c27_r1_io_a),
    .io_s(ft_s5_c27_r1_io_s)
  );
  wire fa_s6_c27_r0_io_a;
  wire fa_s6_c27_r0_io_b;
  wire fa_s6_c27_r0_io_ci;
  wire fa_s6_c27_r0_io_s;
  wire fa_s6_c27_r0_io_co;
  FullAdder fa_s6_c27_r0(
    .io_a(fa_s6_c27_r0_io_a),
    .io_b(fa_s6_c27_r0_io_b),
    .io_ci(fa_s6_c27_r0_io_ci),
    .io_s(fa_s6_c27_r0_io_s),
    .io_co(fa_s6_c27_r0_io_co)
  );
  wire ft_s7_c27_r0_io_a;
  wire ft_s7_c27_r0_io_s;
  FallThrough ft_s7_c27_r0(
    .io_a(ft_s7_c27_r0_io_a),
    .io_s(ft_s7_c27_r0_io_s)
  );
  wire ft_s8_c27_r0_io_a;
  wire ft_s8_c27_r0_io_s;
  FallThrough ft_s8_c27_r0(
    .io_a(ft_s8_c27_r0_io_a),
    .io_s(ft_s8_c27_r0_io_s)
  );
  wire fa_s0_c28_r0_io_a;
  wire fa_s0_c28_r0_io_b;
  wire fa_s0_c28_r0_io_ci;
  wire fa_s0_c28_r0_io_s;
  wire fa_s0_c28_r0_io_co;
  FullAdder fa_s0_c28_r0(
    .io_a(fa_s0_c28_r0_io_a),
    .io_b(fa_s0_c28_r0_io_b),
    .io_ci(fa_s0_c28_r0_io_ci),
    .io_s(fa_s0_c28_r0_io_s),
    .io_co(fa_s0_c28_r0_io_co)
  );
  wire ha_s1_c28_r0_io_a;
  wire ha_s1_c28_r0_io_b;
  wire ha_s1_c28_r0_io_s;
  wire ha_s1_c28_r0_io_co;
  HalfAdder ha_s1_c28_r0(
    .io_a(ha_s1_c28_r0_io_a),
    .io_b(ha_s1_c28_r0_io_b),
    .io_s(ha_s1_c28_r0_io_s),
    .io_co(ha_s1_c28_r0_io_co)
  );
  wire ha_s2_c28_r0_io_a;
  wire ha_s2_c28_r0_io_b;
  wire ha_s2_c28_r0_io_s;
  wire ha_s2_c28_r0_io_co;
  HalfAdder ha_s2_c28_r0(
    .io_a(ha_s2_c28_r0_io_a),
    .io_b(ha_s2_c28_r0_io_b),
    .io_s(ha_s2_c28_r0_io_s),
    .io_co(ha_s2_c28_r0_io_co)
  );
  wire ft_s3_c28_r0_io_a;
  wire ft_s3_c28_r0_io_s;
  FallThrough ft_s3_c28_r0(
    .io_a(ft_s3_c28_r0_io_a),
    .io_s(ft_s3_c28_r0_io_s)
  );
  wire ft_s4_c28_r0_io_a;
  wire ft_s4_c28_r0_io_s;
  FallThrough ft_s4_c28_r0(
    .io_a(ft_s4_c28_r0_io_a),
    .io_s(ft_s4_c28_r0_io_s)
  );
  wire ft_s4_c28_r1_io_a;
  wire ft_s4_c28_r1_io_s;
  FallThrough ft_s4_c28_r1(
    .io_a(ft_s4_c28_r1_io_a),
    .io_s(ft_s4_c28_r1_io_s)
  );
  wire ft_s5_c28_r0_io_a;
  wire ft_s5_c28_r0_io_s;
  FallThrough ft_s5_c28_r0(
    .io_a(ft_s5_c28_r0_io_a),
    .io_s(ft_s5_c28_r0_io_s)
  );
  wire ft_s5_c28_r1_io_a;
  wire ft_s5_c28_r1_io_s;
  FallThrough ft_s5_c28_r1(
    .io_a(ft_s5_c28_r1_io_a),
    .io_s(ft_s5_c28_r1_io_s)
  );
  wire ft_s6_c28_r0_io_a;
  wire ft_s6_c28_r0_io_s;
  FallThrough ft_s6_c28_r0(
    .io_a(ft_s6_c28_r0_io_a),
    .io_s(ft_s6_c28_r0_io_s)
  );
  wire ft_s6_c28_r1_io_a;
  wire ft_s6_c28_r1_io_s;
  FallThrough ft_s6_c28_r1(
    .io_a(ft_s6_c28_r1_io_a),
    .io_s(ft_s6_c28_r1_io_s)
  );
  wire fa_s7_c28_r0_io_a;
  wire fa_s7_c28_r0_io_b;
  wire fa_s7_c28_r0_io_ci;
  wire fa_s7_c28_r0_io_s;
  wire fa_s7_c28_r0_io_co;
  FullAdder fa_s7_c28_r0(
    .io_a(fa_s7_c28_r0_io_a),
    .io_b(fa_s7_c28_r0_io_b),
    .io_ci(fa_s7_c28_r0_io_ci),
    .io_s(fa_s7_c28_r0_io_s),
    .io_co(fa_s7_c28_r0_io_co)
  );
  wire ft_s8_c28_r0_io_a;
  wire ft_s8_c28_r0_io_s;
  FallThrough ft_s8_c28_r0(
    .io_a(ft_s8_c28_r0_io_a),
    .io_s(ft_s8_c28_r0_io_s)
  );
  wire ha_s0_c29_r0_io_a;
  wire ha_s0_c29_r0_io_b;
  wire ha_s0_c29_r0_io_s;
  wire ha_s0_c29_r0_io_co;
  HalfAdder ha_s0_c29_r0(
    .io_a(ha_s0_c29_r0_io_a),
    .io_b(ha_s0_c29_r0_io_b),
    .io_s(ha_s0_c29_r0_io_s),
    .io_co(ha_s0_c29_r0_io_co)
  );
  wire ft_s1_c29_r0_io_a;
  wire ft_s1_c29_r0_io_s;
  FallThrough ft_s1_c29_r0(
    .io_a(ft_s1_c29_r0_io_a),
    .io_s(ft_s1_c29_r0_io_s)
  );
  wire ft_s1_c29_r1_io_a;
  wire ft_s1_c29_r1_io_s;
  FallThrough ft_s1_c29_r1(
    .io_a(ft_s1_c29_r1_io_a),
    .io_s(ft_s1_c29_r1_io_s)
  );
  wire fa_s2_c29_r0_io_a;
  wire fa_s2_c29_r0_io_b;
  wire fa_s2_c29_r0_io_ci;
  wire fa_s2_c29_r0_io_s;
  wire fa_s2_c29_r0_io_co;
  FullAdder fa_s2_c29_r0(
    .io_a(fa_s2_c29_r0_io_a),
    .io_b(fa_s2_c29_r0_io_b),
    .io_ci(fa_s2_c29_r0_io_ci),
    .io_s(fa_s2_c29_r0_io_s),
    .io_co(fa_s2_c29_r0_io_co)
  );
  wire ft_s3_c29_r0_io_a;
  wire ft_s3_c29_r0_io_s;
  FallThrough ft_s3_c29_r0(
    .io_a(ft_s3_c29_r0_io_a),
    .io_s(ft_s3_c29_r0_io_s)
  );
  wire ft_s3_c29_r1_io_a;
  wire ft_s3_c29_r1_io_s;
  FallThrough ft_s3_c29_r1(
    .io_a(ft_s3_c29_r1_io_a),
    .io_s(ft_s3_c29_r1_io_s)
  );
  wire ft_s4_c29_r0_io_a;
  wire ft_s4_c29_r0_io_s;
  FallThrough ft_s4_c29_r0(
    .io_a(ft_s4_c29_r0_io_a),
    .io_s(ft_s4_c29_r0_io_s)
  );
  wire ft_s4_c29_r1_io_a;
  wire ft_s4_c29_r1_io_s;
  FallThrough ft_s4_c29_r1(
    .io_a(ft_s4_c29_r1_io_a),
    .io_s(ft_s4_c29_r1_io_s)
  );
  wire ft_s5_c29_r0_io_a;
  wire ft_s5_c29_r0_io_s;
  FallThrough ft_s5_c29_r0(
    .io_a(ft_s5_c29_r0_io_a),
    .io_s(ft_s5_c29_r0_io_s)
  );
  wire ft_s5_c29_r1_io_a;
  wire ft_s5_c29_r1_io_s;
  FallThrough ft_s5_c29_r1(
    .io_a(ft_s5_c29_r1_io_a),
    .io_s(ft_s5_c29_r1_io_s)
  );
  wire ft_s6_c29_r0_io_a;
  wire ft_s6_c29_r0_io_s;
  FallThrough ft_s6_c29_r0(
    .io_a(ft_s6_c29_r0_io_a),
    .io_s(ft_s6_c29_r0_io_s)
  );
  wire ft_s6_c29_r1_io_a;
  wire ft_s6_c29_r1_io_s;
  FallThrough ft_s6_c29_r1(
    .io_a(ft_s6_c29_r1_io_a),
    .io_s(ft_s6_c29_r1_io_s)
  );
  wire ft_s7_c29_r0_io_a;
  wire ft_s7_c29_r0_io_s;
  FallThrough ft_s7_c29_r0(
    .io_a(ft_s7_c29_r0_io_a),
    .io_s(ft_s7_c29_r0_io_s)
  );
  wire ft_s7_c29_r1_io_a;
  wire ft_s7_c29_r1_io_s;
  FallThrough ft_s7_c29_r1(
    .io_a(ft_s7_c29_r1_io_a),
    .io_s(ft_s7_c29_r1_io_s)
  );
  wire fa_s8_c29_r0_io_a;
  wire fa_s8_c29_r0_io_b;
  wire fa_s8_c29_r0_io_ci;
  wire fa_s8_c29_r0_io_s;
  wire fa_s8_c29_r0_io_co;
  FullAdder fa_s8_c29_r0(
    .io_a(fa_s8_c29_r0_io_a),
    .io_b(fa_s8_c29_r0_io_b),
    .io_ci(fa_s8_c29_r0_io_ci),
    .io_s(fa_s8_c29_r0_io_s),
    .io_co(fa_s8_c29_r0_io_co)
  );
  wire ft_s0_c30_r0_io_a;
  wire ft_s0_c30_r0_io_s;
  FallThrough ft_s0_c30_r0(
    .io_a(ft_s0_c30_r0_io_a),
    .io_s(ft_s0_c30_r0_io_s)
  );
  wire ft_s1_c30_r0_io_a;
  wire ft_s1_c30_r0_io_s;
  FallThrough ft_s1_c30_r0(
    .io_a(ft_s1_c30_r0_io_a),
    .io_s(ft_s1_c30_r0_io_s)
  );
  wire ft_s1_c30_r1_io_a;
  wire ft_s1_c30_r1_io_s;
  FallThrough ft_s1_c30_r1(
    .io_a(ft_s1_c30_r1_io_a),
    .io_s(ft_s1_c30_r1_io_s)
  );
  wire ft_s2_c30_r0_io_a;
  wire ft_s2_c30_r0_io_s;
  FallThrough ft_s2_c30_r0(
    .io_a(ft_s2_c30_r0_io_a),
    .io_s(ft_s2_c30_r0_io_s)
  );
  wire ft_s2_c30_r1_io_a;
  wire ft_s2_c30_r1_io_s;
  FallThrough ft_s2_c30_r1(
    .io_a(ft_s2_c30_r1_io_a),
    .io_s(ft_s2_c30_r1_io_s)
  );
  wire fa_s3_c30_r0_io_a;
  wire fa_s3_c30_r0_io_b;
  wire fa_s3_c30_r0_io_ci;
  wire fa_s3_c30_r0_io_s;
  wire fa_s3_c30_r0_io_co;
  FullAdder fa_s3_c30_r0(
    .io_a(fa_s3_c30_r0_io_a),
    .io_b(fa_s3_c30_r0_io_b),
    .io_ci(fa_s3_c30_r0_io_ci),
    .io_s(fa_s3_c30_r0_io_s),
    .io_co(fa_s3_c30_r0_io_co)
  );
  wire ft_s4_c30_r0_io_a;
  wire ft_s4_c30_r0_io_s;
  FallThrough ft_s4_c30_r0(
    .io_a(ft_s4_c30_r0_io_a),
    .io_s(ft_s4_c30_r0_io_s)
  );
  wire ft_s5_c30_r0_io_a;
  wire ft_s5_c30_r0_io_s;
  FallThrough ft_s5_c30_r0(
    .io_a(ft_s5_c30_r0_io_a),
    .io_s(ft_s5_c30_r0_io_s)
  );
  wire ft_s6_c30_r0_io_a;
  wire ft_s6_c30_r0_io_s;
  FallThrough ft_s6_c30_r0(
    .io_a(ft_s6_c30_r0_io_a),
    .io_s(ft_s6_c30_r0_io_s)
  );
  wire ft_s7_c30_r0_io_a;
  wire ft_s7_c30_r0_io_s;
  FallThrough ft_s7_c30_r0(
    .io_a(ft_s7_c30_r0_io_a),
    .io_s(ft_s7_c30_r0_io_s)
  );
  wire ft_s8_c30_r0_io_a;
  wire ft_s8_c30_r0_io_s;
  FallThrough ft_s8_c30_r0(
    .io_a(ft_s8_c30_r0_io_a),
    .io_s(ft_s8_c30_r0_io_s)
  );
  wire ft_s4_c31_r0_io_a;
  wire ft_s4_c31_r0_io_s;
  FallThrough ft_s4_c31_r0(
    .io_a(ft_s4_c31_r0_io_a),
    .io_s(ft_s4_c31_r0_io_s)
  );
  wire ft_s5_c31_r0_io_a;
  wire ft_s5_c31_r0_io_s;
  FallThrough ft_s5_c31_r0(
    .io_a(ft_s5_c31_r0_io_a),
    .io_s(ft_s5_c31_r0_io_s)
  );
  wire ft_s6_c31_r0_io_a;
  wire ft_s6_c31_r0_io_s;
  FallThrough ft_s6_c31_r0(
    .io_a(ft_s6_c31_r0_io_a),
    .io_s(ft_s6_c31_r0_io_s)
  );
  wire ft_s7_c31_r0_io_a;
  wire ft_s7_c31_r0_io_s;
  FallThrough ft_s7_c31_r0(
    .io_a(ft_s7_c31_r0_io_a),
    .io_s(ft_s7_c31_r0_io_s)
  );
  wire ft_s8_c31_r0_io_a;
  wire ft_s8_c31_r0_io_s;
  FallThrough ft_s8_c31_r0(
    .io_a(ft_s8_c31_r0_io_a),
    .io_s(ft_s8_c31_r0_io_s)
  );
  assign ft_s0_c0_r0_io_a = io_pp_0[0];
  assign ha_s0_c1_r0_io_a = io_pp_1[0];
  assign ha_s0_c1_r0_io_b = io_pp_1[1];
  assign ha_s0_c2_r0_io_a = io_pp_2[0];
  assign ha_s0_c2_r0_io_b = io_pp_2[1];
  assign ft_s0_c2_r1_io_a = io_pp_2[2];
  assign fa_s0_c3_r0_io_a = io_pp_3[0];
  assign fa_s0_c3_r0_io_b = io_pp_3[1];
  assign fa_s0_c3_r0_io_ci = io_pp_3[2];
  assign ft_s0_c3_r1_io_a = io_pp_3[3];
  assign fa_s0_c4_r0_io_a = io_pp_4[0];
  assign fa_s0_c4_r0_io_b = io_pp_4[1];
  assign fa_s0_c4_r0_io_ci = io_pp_4[2];
  assign ft_s0_c4_r1_io_a = io_pp_4[3];
  assign ft_s0_c4_r2_io_a = io_pp_4[4];
  assign fa_s0_c5_r0_io_a = io_pp_5[0];
  assign fa_s0_c5_r0_io_b = io_pp_5[1];
  assign fa_s0_c5_r0_io_ci = io_pp_5[2];
  assign fa_s0_c5_r1_io_a = io_pp_5[3];
  assign fa_s0_c5_r1_io_b = io_pp_5[4];
  assign fa_s0_c5_r1_io_ci = io_pp_5[5];
  assign fa_s0_c6_r0_io_a = io_pp_6[0];
  assign fa_s0_c6_r0_io_b = io_pp_6[1];
  assign fa_s0_c6_r0_io_ci = io_pp_6[2];
  assign fa_s0_c6_r1_io_a = io_pp_6[3];
  assign fa_s0_c6_r1_io_b = io_pp_6[4];
  assign fa_s0_c6_r1_io_ci = io_pp_6[5];
  assign ft_s0_c6_r2_io_a = io_pp_6[6];
  assign fa_s0_c7_r0_io_a = io_pp_7[0];
  assign fa_s0_c7_r0_io_b = io_pp_7[1];
  assign fa_s0_c7_r0_io_ci = io_pp_7[2];
  assign fa_s0_c7_r1_io_a = io_pp_7[3];
  assign fa_s0_c7_r1_io_b = io_pp_7[4];
  assign fa_s0_c7_r1_io_ci = io_pp_7[5];
  assign ft_s0_c7_r2_io_a = io_pp_7[6];
  assign ft_s0_c7_r3_io_a = io_pp_7[7];
  assign fa_s0_c8_r0_io_a = io_pp_8[0];
  assign fa_s0_c8_r0_io_b = io_pp_8[1];
  assign fa_s0_c8_r0_io_ci = io_pp_8[2];
  assign fa_s0_c8_r1_io_a = io_pp_8[3];
  assign fa_s0_c8_r1_io_b = io_pp_8[4];
  assign fa_s0_c8_r1_io_ci = io_pp_8[5];
  assign fa_s0_c8_r2_io_a = io_pp_8[6];
  assign fa_s0_c8_r2_io_b = io_pp_8[7];
  assign fa_s0_c8_r2_io_ci = io_pp_8[8];
  assign fa_s0_c9_r0_io_a = io_pp_9[0];
  assign fa_s0_c9_r0_io_b = io_pp_9[1];
  assign fa_s0_c9_r0_io_ci = io_pp_9[2];
  assign fa_s0_c9_r1_io_a = io_pp_9[3];
  assign fa_s0_c9_r1_io_b = io_pp_9[4];
  assign fa_s0_c9_r1_io_ci = io_pp_9[5];
  assign fa_s0_c9_r2_io_a = io_pp_9[6];
  assign fa_s0_c9_r2_io_b = io_pp_9[7];
  assign fa_s0_c9_r2_io_ci = io_pp_9[8];
  assign ft_s0_c9_r3_io_a = io_pp_9[9];
  assign fa_s0_c10_r0_io_a = io_pp_10[0];
  assign fa_s0_c10_r0_io_b = io_pp_10[1];
  assign fa_s0_c10_r0_io_ci = io_pp_10[2];
  assign fa_s0_c10_r1_io_a = io_pp_10[3];
  assign fa_s0_c10_r1_io_b = io_pp_10[4];
  assign fa_s0_c10_r1_io_ci = io_pp_10[5];
  assign fa_s0_c10_r2_io_a = io_pp_10[6];
  assign fa_s0_c10_r2_io_b = io_pp_10[7];
  assign fa_s0_c10_r2_io_ci = io_pp_10[8];
  assign ft_s0_c10_r3_io_a = io_pp_10[9];
  assign ft_s0_c10_r4_io_a = io_pp_10[10];
  assign fa_s0_c11_r0_io_a = io_pp_11[0];
  assign fa_s0_c11_r0_io_b = io_pp_11[1];
  assign fa_s0_c11_r0_io_ci = io_pp_11[2];
  assign fa_s0_c11_r1_io_a = io_pp_11[3];
  assign fa_s0_c11_r1_io_b = io_pp_11[4];
  assign fa_s0_c11_r1_io_ci = io_pp_11[5];
  assign fa_s0_c11_r2_io_a = io_pp_11[6];
  assign fa_s0_c11_r2_io_b = io_pp_11[7];
  assign fa_s0_c11_r2_io_ci = io_pp_11[8];
  assign fa_s0_c11_r3_io_a = io_pp_11[9];
  assign fa_s0_c11_r3_io_b = io_pp_11[10];
  assign fa_s0_c11_r3_io_ci = io_pp_11[11];
  assign fa_s0_c12_r0_io_a = io_pp_12[0];
  assign fa_s0_c12_r0_io_b = io_pp_12[1];
  assign fa_s0_c12_r0_io_ci = io_pp_12[2];
  assign fa_s0_c12_r1_io_a = io_pp_12[3];
  assign fa_s0_c12_r1_io_b = io_pp_12[4];
  assign fa_s0_c12_r1_io_ci = io_pp_12[5];
  assign fa_s0_c12_r2_io_a = io_pp_12[6];
  assign fa_s0_c12_r2_io_b = io_pp_12[7];
  assign fa_s0_c12_r2_io_ci = io_pp_12[8];
  assign fa_s0_c12_r3_io_a = io_pp_12[9];
  assign fa_s0_c12_r3_io_b = io_pp_12[10];
  assign fa_s0_c12_r3_io_ci = io_pp_12[11];
  assign ft_s0_c12_r4_io_a = io_pp_12[12];
  assign fa_s0_c13_r0_io_a = io_pp_13[0];
  assign fa_s0_c13_r0_io_b = io_pp_13[1];
  assign fa_s0_c13_r0_io_ci = io_pp_13[2];
  assign fa_s0_c13_r1_io_a = io_pp_13[3];
  assign fa_s0_c13_r1_io_b = io_pp_13[4];
  assign fa_s0_c13_r1_io_ci = io_pp_13[5];
  assign fa_s0_c13_r2_io_a = io_pp_13[6];
  assign fa_s0_c13_r2_io_b = io_pp_13[7];
  assign fa_s0_c13_r2_io_ci = io_pp_13[8];
  assign fa_s0_c13_r3_io_a = io_pp_13[9];
  assign fa_s0_c13_r3_io_b = io_pp_13[10];
  assign fa_s0_c13_r3_io_ci = io_pp_13[11];
  assign ft_s0_c13_r4_io_a = io_pp_13[12];
  assign ft_s0_c13_r5_io_a = io_pp_13[13];
  assign fa_s0_c14_r0_io_a = io_pp_14[0];
  assign fa_s0_c14_r0_io_b = io_pp_14[1];
  assign fa_s0_c14_r0_io_ci = io_pp_14[2];
  assign fa_s0_c14_r1_io_a = io_pp_14[3];
  assign fa_s0_c14_r1_io_b = io_pp_14[4];
  assign fa_s0_c14_r1_io_ci = io_pp_14[5];
  assign fa_s0_c14_r2_io_a = io_pp_14[6];
  assign fa_s0_c14_r2_io_b = io_pp_14[7];
  assign fa_s0_c14_r2_io_ci = io_pp_14[8];
  assign fa_s0_c14_r3_io_a = io_pp_14[9];
  assign fa_s0_c14_r3_io_b = io_pp_14[10];
  assign fa_s0_c14_r3_io_ci = io_pp_14[11];
  assign fa_s0_c14_r4_io_a = io_pp_14[12];
  assign fa_s0_c14_r4_io_b = io_pp_14[13];
  assign fa_s0_c14_r4_io_ci = io_pp_14[14];
  assign fa_s0_c15_r0_io_a = io_pp_15[0];
  assign fa_s0_c15_r0_io_b = io_pp_15[1];
  assign fa_s0_c15_r0_io_ci = io_pp_15[2];
  assign fa_s0_c15_r1_io_a = io_pp_15[3];
  assign fa_s0_c15_r1_io_b = io_pp_15[4];
  assign fa_s0_c15_r1_io_ci = io_pp_15[5];
  assign fa_s0_c15_r2_io_a = io_pp_15[6];
  assign fa_s0_c15_r2_io_b = io_pp_15[7];
  assign fa_s0_c15_r2_io_ci = io_pp_15[8];
  assign fa_s0_c15_r3_io_a = io_pp_15[9];
  assign fa_s0_c15_r3_io_b = io_pp_15[10];
  assign fa_s0_c15_r3_io_ci = io_pp_15[11];
  assign fa_s0_c15_r4_io_a = io_pp_15[12];
  assign fa_s0_c15_r4_io_b = io_pp_15[13];
  assign fa_s0_c15_r4_io_ci = io_pp_15[14];
  assign ft_s0_c15_r5_io_a = io_pp_15[15];
  assign fa_s0_c16_r0_io_a = io_pp_16[0];
  assign fa_s0_c16_r0_io_b = io_pp_16[1];
  assign fa_s0_c16_r0_io_ci = io_pp_16[2];
  assign fa_s0_c16_r1_io_a = io_pp_16[3];
  assign fa_s0_c16_r1_io_b = io_pp_16[4];
  assign fa_s0_c16_r1_io_ci = io_pp_16[5];
  assign fa_s0_c16_r2_io_a = io_pp_16[6];
  assign fa_s0_c16_r2_io_b = io_pp_16[7];
  assign fa_s0_c16_r2_io_ci = io_pp_16[8];
  assign fa_s0_c16_r3_io_a = io_pp_16[9];
  assign fa_s0_c16_r3_io_b = io_pp_16[10];
  assign fa_s0_c16_r3_io_ci = io_pp_16[11];
  assign fa_s0_c16_r4_io_a = io_pp_16[12];
  assign fa_s0_c16_r4_io_b = io_pp_16[13];
  assign fa_s0_c16_r4_io_ci = io_pp_16[14];
  assign fa_s0_c17_r0_io_a = io_pp_17[0];
  assign fa_s0_c17_r0_io_b = io_pp_17[1];
  assign fa_s0_c17_r0_io_ci = io_pp_17[2];
  assign fa_s0_c17_r1_io_a = io_pp_17[3];
  assign fa_s0_c17_r1_io_b = io_pp_17[4];
  assign fa_s0_c17_r1_io_ci = io_pp_17[5];
  assign fa_s0_c17_r2_io_a = io_pp_17[6];
  assign fa_s0_c17_r2_io_b = io_pp_17[7];
  assign fa_s0_c17_r2_io_ci = io_pp_17[8];
  assign fa_s0_c17_r3_io_a = io_pp_17[9];
  assign fa_s0_c17_r3_io_b = io_pp_17[10];
  assign fa_s0_c17_r3_io_ci = io_pp_17[11];
  assign ft_s0_c17_r4_io_a = io_pp_17[12];
  assign ft_s0_c17_r5_io_a = io_pp_17[13];
  assign fa_s0_c18_r0_io_a = io_pp_18[0];
  assign fa_s0_c18_r0_io_b = io_pp_18[1];
  assign fa_s0_c18_r0_io_ci = io_pp_18[2];
  assign fa_s0_c18_r1_io_a = io_pp_18[3];
  assign fa_s0_c18_r1_io_b = io_pp_18[4];
  assign fa_s0_c18_r1_io_ci = io_pp_18[5];
  assign fa_s0_c18_r2_io_a = io_pp_18[6];
  assign fa_s0_c18_r2_io_b = io_pp_18[7];
  assign fa_s0_c18_r2_io_ci = io_pp_18[8];
  assign fa_s0_c18_r3_io_a = io_pp_18[9];
  assign fa_s0_c18_r3_io_b = io_pp_18[10];
  assign fa_s0_c18_r3_io_ci = io_pp_18[11];
  assign ft_s0_c18_r4_io_a = io_pp_18[12];
  assign fa_s0_c19_r0_io_a = io_pp_19[0];
  assign fa_s0_c19_r0_io_b = io_pp_19[1];
  assign fa_s0_c19_r0_io_ci = io_pp_19[2];
  assign fa_s0_c19_r1_io_a = io_pp_19[3];
  assign fa_s0_c19_r1_io_b = io_pp_19[4];
  assign fa_s0_c19_r1_io_ci = io_pp_19[5];
  assign fa_s0_c19_r2_io_a = io_pp_19[6];
  assign fa_s0_c19_r2_io_b = io_pp_19[7];
  assign fa_s0_c19_r2_io_ci = io_pp_19[8];
  assign fa_s0_c19_r3_io_a = io_pp_19[9];
  assign fa_s0_c19_r3_io_b = io_pp_19[10];
  assign fa_s0_c19_r3_io_ci = io_pp_19[11];
  assign fa_s0_c20_r0_io_a = io_pp_20[0];
  assign fa_s0_c20_r0_io_b = io_pp_20[1];
  assign fa_s0_c20_r0_io_ci = io_pp_20[2];
  assign fa_s0_c20_r1_io_a = io_pp_20[3];
  assign fa_s0_c20_r1_io_b = io_pp_20[4];
  assign fa_s0_c20_r1_io_ci = io_pp_20[5];
  assign fa_s0_c20_r2_io_a = io_pp_20[6];
  assign fa_s0_c20_r2_io_b = io_pp_20[7];
  assign fa_s0_c20_r2_io_ci = io_pp_20[8];
  assign ha_s0_c20_r3_io_a = io_pp_20[9];
  assign ha_s0_c20_r3_io_b = io_pp_20[10];
  assign fa_s0_c21_r0_io_a = io_pp_21[0];
  assign fa_s0_c21_r0_io_b = io_pp_21[1];
  assign fa_s0_c21_r0_io_ci = io_pp_21[2];
  assign fa_s0_c21_r1_io_a = io_pp_21[3];
  assign fa_s0_c21_r1_io_b = io_pp_21[4];
  assign fa_s0_c21_r1_io_ci = io_pp_21[5];
  assign fa_s0_c21_r2_io_a = io_pp_21[6];
  assign fa_s0_c21_r2_io_b = io_pp_21[7];
  assign fa_s0_c21_r2_io_ci = io_pp_21[8];
  assign ft_s0_c21_r3_io_a = io_pp_21[9];
  assign fa_s0_c22_r0_io_a = io_pp_22[0];
  assign fa_s0_c22_r0_io_b = io_pp_22[1];
  assign fa_s0_c22_r0_io_ci = io_pp_22[2];
  assign fa_s0_c22_r1_io_a = io_pp_22[3];
  assign fa_s0_c22_r1_io_b = io_pp_22[4];
  assign fa_s0_c22_r1_io_ci = io_pp_22[5];
  assign fa_s0_c22_r2_io_a = io_pp_22[6];
  assign fa_s0_c22_r2_io_b = io_pp_22[7];
  assign fa_s0_c22_r2_io_ci = io_pp_22[8];
  assign fa_s0_c23_r0_io_a = io_pp_23[0];
  assign fa_s0_c23_r0_io_b = io_pp_23[1];
  assign fa_s0_c23_r0_io_ci = io_pp_23[2];
  assign fa_s0_c23_r1_io_a = io_pp_23[3];
  assign fa_s0_c23_r1_io_b = io_pp_23[4];
  assign fa_s0_c23_r1_io_ci = io_pp_23[5];
  assign ft_s0_c23_r2_io_a = io_pp_23[6];
  assign ft_s0_c23_r3_io_a = io_pp_23[7];
  assign fa_s0_c24_r0_io_a = io_pp_24[0];
  assign fa_s0_c24_r0_io_b = io_pp_24[1];
  assign fa_s0_c24_r0_io_ci = io_pp_24[2];
  assign fa_s0_c24_r1_io_a = io_pp_24[3];
  assign fa_s0_c24_r1_io_b = io_pp_24[4];
  assign fa_s0_c24_r1_io_ci = io_pp_24[5];
  assign ft_s0_c24_r2_io_a = io_pp_24[6];
  assign fa_s0_c25_r0_io_a = io_pp_25[0];
  assign fa_s0_c25_r0_io_b = io_pp_25[1];
  assign fa_s0_c25_r0_io_ci = io_pp_25[2];
  assign fa_s0_c25_r1_io_a = io_pp_25[3];
  assign fa_s0_c25_r1_io_b = io_pp_25[4];
  assign fa_s0_c25_r1_io_ci = io_pp_25[5];
  assign fa_s0_c26_r0_io_a = io_pp_26[0];
  assign fa_s0_c26_r0_io_b = io_pp_26[1];
  assign fa_s0_c26_r0_io_ci = io_pp_26[2];
  assign ft_s0_c26_r1_io_a = io_pp_26[3];
  assign ft_s0_c26_r2_io_a = io_pp_26[4];
  assign fa_s0_c27_r0_io_a = io_pp_27[0];
  assign fa_s0_c27_r0_io_b = io_pp_27[1];
  assign fa_s0_c27_r0_io_ci = io_pp_27[2];
  assign ft_s0_c27_r1_io_a = io_pp_27[3];
  assign fa_s0_c28_r0_io_a = io_pp_28[0];
  assign fa_s0_c28_r0_io_b = io_pp_28[1];
  assign fa_s0_c28_r0_io_ci = io_pp_28[2];
  assign ha_s0_c29_r0_io_a = io_pp_29[0];
  assign ha_s0_c29_r0_io_b = io_pp_29[1];
  assign ft_s0_c30_r0_io_a = io_pp_30[0];
  assign ft_s1_c0_r0_io_a = ft_s0_c0_r0_io_s;
  assign ft_s2_c0_r0_io_a = ft_s1_c0_r0_io_s;
  assign ft_s3_c0_r0_io_a = ft_s2_c0_r0_io_s;
  assign ft_s4_c0_r0_io_a = ft_s3_c0_r0_io_s;
  assign ft_s5_c0_r0_io_a = ft_s4_c0_r0_io_s;
  assign ft_s6_c0_r0_io_a = ft_s5_c0_r0_io_s;
  assign ft_s7_c0_r0_io_a = ft_s6_c0_r0_io_s;
  assign ft_s8_c0_r0_io_a = ft_s7_c0_r0_io_s;
  assign io_augend[0] = ft_s8_c0_r0_io_s;
  assign ft_s1_c1_r0_io_a = ha_s0_c1_r0_io_s;
  assign ft_s1_c2_r1_io_a = ha_s0_c1_r0_io_co;
  assign ft_s2_c1_r0_io_a = ft_s1_c1_r0_io_s;
  assign ft_s3_c1_r0_io_a = ft_s2_c1_r0_io_s;
  assign ft_s4_c1_r0_io_a = ft_s3_c1_r0_io_s;
  assign ft_s5_c1_r0_io_a = ft_s4_c1_r0_io_s;
  assign ft_s6_c1_r0_io_a = ft_s5_c1_r0_io_s;
  assign ft_s7_c1_r0_io_a = ft_s6_c1_r0_io_s;
  assign ft_s8_c1_r0_io_a = ft_s7_c1_r0_io_s;
  assign io_augend[1] = ft_s8_c1_r0_io_s;
  assign ha_s1_c2_r0_io_a = ha_s0_c2_r0_io_s;
  assign fa_s1_c3_r0_io_ci = ha_s0_c2_r0_io_co;
  assign ha_s1_c2_r0_io_b = ft_s0_c2_r1_io_s;
  assign ft_s2_c2_r0_io_a = ha_s1_c2_r0_io_s;
  assign ha_s2_c3_r0_io_b = ha_s1_c2_r0_io_co;
  assign ft_s2_c2_r1_io_a = ft_s1_c2_r1_io_s;
  assign ft_s3_c2_r0_io_a = ft_s2_c2_r0_io_s;
  assign ft_s3_c2_r1_io_a = ft_s2_c2_r1_io_s;
  assign ft_s4_c2_r0_io_a = ft_s3_c2_r0_io_s;
  assign ft_s4_c2_r1_io_a = ft_s3_c2_r1_io_s;
  assign ft_s5_c2_r0_io_a = ft_s4_c2_r0_io_s;
  assign ft_s5_c2_r1_io_a = ft_s4_c2_r1_io_s;
  assign ft_s6_c2_r0_io_a = ft_s5_c2_r0_io_s;
  assign ft_s6_c2_r1_io_a = ft_s5_c2_r1_io_s;
  assign ft_s7_c2_r0_io_a = ft_s6_c2_r0_io_s;
  assign ft_s7_c2_r1_io_a = ft_s6_c2_r1_io_s;
  assign ft_s8_c2_r0_io_a = ft_s7_c2_r0_io_s;
  assign ft_s8_c2_r1_io_a = ft_s7_c2_r1_io_s;
  assign io_augend[2] = ft_s8_c2_r0_io_s;
  assign io_addend[2] = ft_s8_c2_r1_io_s;
  assign fa_s1_c3_r0_io_a = fa_s0_c3_r0_io_s;
  assign ft_s1_c4_r1_io_a = fa_s0_c3_r0_io_co;
  assign fa_s1_c3_r0_io_b = ft_s0_c3_r1_io_s;
  assign ha_s2_c3_r0_io_a = fa_s1_c3_r0_io_s;
  assign fa_s2_c4_r0_io_ci = fa_s1_c3_r0_io_co;
  assign ft_s3_c3_r0_io_a = ha_s2_c3_r0_io_s;
  assign ft_s3_c4_r1_io_a = ha_s2_c3_r0_io_co;
  assign ft_s4_c3_r0_io_a = ft_s3_c3_r0_io_s;
  assign ft_s5_c3_r0_io_a = ft_s4_c3_r0_io_s;
  assign ft_s6_c3_r0_io_a = ft_s5_c3_r0_io_s;
  assign ft_s7_c3_r0_io_a = ft_s6_c3_r0_io_s;
  assign ft_s8_c3_r0_io_a = ft_s7_c3_r0_io_s;
  assign io_augend[3] = ft_s8_c3_r0_io_s;
  assign fa_s1_c4_r0_io_a = fa_s0_c4_r0_io_s;
  assign fa_s1_c5_r0_io_ci = fa_s0_c4_r0_io_co;
  assign fa_s1_c4_r0_io_b = ft_s0_c4_r1_io_s;
  assign fa_s1_c4_r0_io_ci = ft_s0_c4_r2_io_s;
  assign fa_s2_c4_r0_io_a = fa_s1_c4_r0_io_s;
  assign ft_s2_c5_r1_io_a = fa_s1_c4_r0_io_co;
  assign fa_s2_c4_r0_io_b = ft_s1_c4_r1_io_s;
  assign ft_s3_c4_r0_io_a = fa_s2_c4_r0_io_s;
  assign fa_s3_c5_r0_io_ci = fa_s2_c4_r0_io_co;
  assign ft_s4_c4_r0_io_a = ft_s3_c4_r0_io_s;
  assign ft_s4_c4_r1_io_a = ft_s3_c4_r1_io_s;
  assign ft_s5_c4_r0_io_a = ft_s4_c4_r0_io_s;
  assign ft_s5_c4_r1_io_a = ft_s4_c4_r1_io_s;
  assign ft_s6_c4_r0_io_a = ft_s5_c4_r0_io_s;
  assign ft_s6_c4_r1_io_a = ft_s5_c4_r1_io_s;
  assign ft_s7_c4_r0_io_a = ft_s6_c4_r0_io_s;
  assign ft_s7_c4_r1_io_a = ft_s6_c4_r1_io_s;
  assign ft_s8_c4_r0_io_a = ft_s7_c4_r0_io_s;
  assign ft_s8_c4_r1_io_a = ft_s7_c4_r1_io_s;
  assign io_augend[4] = ft_s8_c4_r0_io_s;
  assign io_addend[4] = ft_s8_c4_r1_io_s;
  assign fa_s1_c5_r0_io_a = fa_s0_c5_r0_io_s;
  assign ha_s1_c6_r1_io_a = fa_s0_c5_r0_io_co;
  assign fa_s1_c5_r0_io_b = fa_s0_c5_r1_io_s;
  assign ha_s1_c6_r1_io_b = fa_s0_c5_r1_io_co;
  assign ft_s2_c5_r0_io_a = fa_s1_c5_r0_io_s;
  assign fa_s2_c6_r0_io_ci = fa_s1_c5_r0_io_co;
  assign fa_s3_c5_r0_io_a = ft_s2_c5_r0_io_s;
  assign fa_s3_c5_r0_io_b = ft_s2_c5_r1_io_s;
  assign ft_s4_c5_r0_io_a = fa_s3_c5_r0_io_s;
  assign ft_s4_c6_r1_io_a = fa_s3_c5_r0_io_co;
  assign ft_s5_c5_r0_io_a = ft_s4_c5_r0_io_s;
  assign ft_s6_c5_r0_io_a = ft_s5_c5_r0_io_s;
  assign ft_s7_c5_r0_io_a = ft_s6_c5_r0_io_s;
  assign ft_s8_c5_r0_io_a = ft_s7_c5_r0_io_s;
  assign io_augend[5] = ft_s8_c5_r0_io_s;
  assign fa_s1_c6_r0_io_a = fa_s0_c6_r0_io_s;
  assign fa_s1_c7_r1_io_b = fa_s0_c6_r0_io_co;
  assign fa_s1_c6_r0_io_b = fa_s0_c6_r1_io_s;
  assign fa_s1_c7_r1_io_ci = fa_s0_c6_r1_io_co;
  assign fa_s1_c6_r0_io_ci = ft_s0_c6_r2_io_s;
  assign fa_s2_c6_r0_io_a = fa_s1_c6_r0_io_s;
  assign fa_s2_c7_r0_io_ci = fa_s1_c6_r0_io_co;
  assign fa_s2_c6_r0_io_b = ha_s1_c6_r1_io_s;
  assign ft_s2_c7_r1_io_a = ha_s1_c6_r1_io_co;
  assign ft_s3_c6_r0_io_a = fa_s2_c6_r0_io_s;
  assign fa_s3_c7_r0_io_ci = fa_s2_c6_r0_io_co;
  assign ft_s4_c6_r0_io_a = ft_s3_c6_r0_io_s;
  assign ft_s5_c6_r0_io_a = ft_s4_c6_r0_io_s;
  assign ft_s5_c6_r1_io_a = ft_s4_c6_r1_io_s;
  assign ft_s6_c6_r0_io_a = ft_s5_c6_r0_io_s;
  assign ft_s6_c6_r1_io_a = ft_s5_c6_r1_io_s;
  assign ft_s7_c6_r0_io_a = ft_s6_c6_r0_io_s;
  assign ft_s7_c6_r1_io_a = ft_s6_c6_r1_io_s;
  assign ft_s8_c6_r0_io_a = ft_s7_c6_r0_io_s;
  assign ft_s8_c6_r1_io_a = ft_s7_c6_r1_io_s;
  assign io_augend[6] = ft_s8_c6_r0_io_s;
  assign io_addend[6] = ft_s8_c6_r1_io_s;
  assign fa_s1_c7_r0_io_a = fa_s0_c7_r0_io_s;
  assign ha_s1_c8_r1_io_a = fa_s0_c7_r0_io_co;
  assign fa_s1_c7_r0_io_b = fa_s0_c7_r1_io_s;
  assign ha_s1_c8_r1_io_b = fa_s0_c7_r1_io_co;
  assign fa_s1_c7_r0_io_ci = ft_s0_c7_r2_io_s;
  assign fa_s1_c7_r1_io_a = ft_s0_c7_r3_io_s;
  assign fa_s2_c7_r0_io_a = fa_s1_c7_r0_io_s;
  assign fa_s2_c8_r0_io_ci = fa_s1_c7_r0_io_co;
  assign fa_s2_c7_r0_io_b = fa_s1_c7_r1_io_s;
  assign ft_s2_c8_r1_io_a = fa_s1_c7_r1_io_co;
  assign fa_s3_c7_r0_io_a = fa_s2_c7_r0_io_s;
  assign fa_s3_c8_r0_io_ci = fa_s2_c7_r0_io_co;
  assign fa_s3_c7_r0_io_b = ft_s2_c7_r1_io_s;
  assign ft_s4_c7_r0_io_a = fa_s3_c7_r0_io_s;
  assign ft_s4_c8_r1_io_a = fa_s3_c7_r0_io_co;
  assign ft_s5_c7_r0_io_a = ft_s4_c7_r0_io_s;
  assign ft_s6_c7_r0_io_a = ft_s5_c7_r0_io_s;
  assign ft_s7_c7_r0_io_a = ft_s6_c7_r0_io_s;
  assign ft_s8_c7_r0_io_a = ft_s7_c7_r0_io_s;
  assign io_augend[7] = ft_s8_c7_r0_io_s;
  assign fa_s1_c8_r0_io_a = fa_s0_c8_r0_io_s;
  assign fa_s1_c9_r1_io_b = fa_s0_c8_r0_io_co;
  assign fa_s1_c8_r0_io_b = fa_s0_c8_r1_io_s;
  assign fa_s1_c9_r1_io_ci = fa_s0_c8_r1_io_co;
  assign fa_s1_c8_r0_io_ci = fa_s0_c8_r2_io_s;
  assign ft_s1_c9_r2_io_a = fa_s0_c8_r2_io_co;
  assign fa_s2_c8_r0_io_a = fa_s1_c8_r0_io_s;
  assign ha_s2_c9_r1_io_b = fa_s1_c8_r0_io_co;
  assign fa_s2_c8_r0_io_b = ha_s1_c8_r1_io_s;
  assign ft_s2_c9_r2_io_a = ha_s1_c8_r1_io_co;
  assign fa_s3_c8_r0_io_a = fa_s2_c8_r0_io_s;
  assign ft_s3_c9_r2_io_a = fa_s2_c8_r0_io_co;
  assign fa_s3_c8_r0_io_b = ft_s2_c8_r1_io_s;
  assign ft_s4_c8_r0_io_a = fa_s3_c8_r0_io_s;
  assign ft_s4_c9_r2_io_a = fa_s3_c8_r0_io_co;
  assign ft_s5_c8_r0_io_a = ft_s4_c8_r0_io_s;
  assign ft_s5_c8_r1_io_a = ft_s4_c8_r1_io_s;
  assign ft_s6_c8_r0_io_a = ft_s5_c8_r0_io_s;
  assign ft_s6_c8_r1_io_a = ft_s5_c8_r1_io_s;
  assign ft_s7_c8_r0_io_a = ft_s6_c8_r0_io_s;
  assign ft_s7_c8_r1_io_a = ft_s6_c8_r1_io_s;
  assign ft_s8_c8_r0_io_a = ft_s7_c8_r0_io_s;
  assign ft_s8_c8_r1_io_a = ft_s7_c8_r1_io_s;
  assign io_augend[8] = ft_s8_c8_r0_io_s;
  assign io_addend[8] = ft_s8_c8_r1_io_s;
  assign fa_s1_c9_r0_io_a = fa_s0_c9_r0_io_s;
  assign fa_s1_c10_r1_io_ci = fa_s0_c9_r0_io_co;
  assign fa_s1_c9_r0_io_b = fa_s0_c9_r1_io_s;
  assign ft_s1_c10_r2_io_a = fa_s0_c9_r1_io_co;
  assign fa_s1_c9_r0_io_ci = fa_s0_c9_r2_io_s;
  assign ft_s1_c10_r3_io_a = fa_s0_c9_r2_io_co;
  assign fa_s1_c9_r1_io_a = ft_s0_c9_r3_io_s;
  assign ha_s2_c9_r0_io_a = fa_s1_c9_r0_io_s;
  assign fa_s2_c10_r1_io_b = fa_s1_c9_r0_io_co;
  assign ha_s2_c9_r0_io_b = fa_s1_c9_r1_io_s;
  assign fa_s2_c10_r1_io_ci = fa_s1_c9_r1_io_co;
  assign ha_s2_c9_r1_io_a = ft_s1_c9_r2_io_s;
  assign ha_s3_c9_r0_io_a = ha_s2_c9_r0_io_s;
  assign fa_s3_c10_r0_io_ci = ha_s2_c9_r0_io_co;
  assign ha_s3_c9_r0_io_b = ha_s2_c9_r1_io_s;
  assign ft_s3_c10_r1_io_a = ha_s2_c9_r1_io_co;
  assign ft_s3_c9_r1_io_a = ft_s2_c9_r2_io_s;
  assign ha_s4_c9_r0_io_a = ha_s3_c9_r0_io_s;
  assign fa_s4_c10_r0_io_ci = ha_s3_c9_r0_io_co;
  assign ha_s4_c9_r0_io_b = ft_s3_c9_r1_io_s;
  assign ft_s4_c9_r1_io_a = ft_s3_c9_r2_io_s;
  assign fa_s5_c9_r0_io_a = ha_s4_c9_r0_io_s;
  assign ft_s5_c10_r1_io_a = ha_s4_c9_r0_io_co;
  assign fa_s5_c9_r0_io_b = ft_s4_c9_r1_io_s;
  assign fa_s5_c9_r0_io_ci = ft_s4_c9_r2_io_s;
  assign ft_s6_c9_r0_io_a = fa_s5_c9_r0_io_s;
  assign fa_s6_c10_r0_io_ci = fa_s5_c9_r0_io_co;
  assign ft_s7_c9_r0_io_a = ft_s6_c9_r0_io_s;
  assign ft_s8_c9_r0_io_a = ft_s7_c9_r0_io_s;
  assign io_augend[9] = ft_s8_c9_r0_io_s;
  assign fa_s1_c10_r0_io_a = fa_s0_c10_r0_io_s;
  assign fa_s1_c11_r1_io_b = fa_s0_c10_r0_io_co;
  assign fa_s1_c10_r0_io_b = fa_s0_c10_r1_io_s;
  assign fa_s1_c11_r1_io_ci = fa_s0_c10_r1_io_co;
  assign fa_s1_c10_r0_io_ci = fa_s0_c10_r2_io_s;
  assign ft_s1_c11_r2_io_a = fa_s0_c10_r2_io_co;
  assign fa_s1_c10_r1_io_a = ft_s0_c10_r3_io_s;
  assign fa_s1_c10_r1_io_b = ft_s0_c10_r4_io_s;
  assign fa_s2_c10_r0_io_a = fa_s1_c10_r0_io_s;
  assign ha_s2_c11_r1_io_a = fa_s1_c10_r0_io_co;
  assign fa_s2_c10_r0_io_b = fa_s1_c10_r1_io_s;
  assign ha_s2_c11_r1_io_b = fa_s1_c10_r1_io_co;
  assign fa_s2_c10_r0_io_ci = ft_s1_c10_r2_io_s;
  assign fa_s2_c10_r1_io_a = ft_s1_c10_r3_io_s;
  assign fa_s3_c10_r0_io_a = fa_s2_c10_r0_io_s;
  assign fa_s3_c11_r0_io_ci = fa_s2_c10_r0_io_co;
  assign fa_s3_c10_r0_io_b = fa_s2_c10_r1_io_s;
  assign ft_s3_c11_r1_io_a = fa_s2_c10_r1_io_co;
  assign fa_s4_c10_r0_io_a = fa_s3_c10_r0_io_s;
  assign ft_s4_c11_r1_io_a = fa_s3_c10_r0_io_co;
  assign fa_s4_c10_r0_io_b = ft_s3_c10_r1_io_s;
  assign ft_s5_c10_r0_io_a = fa_s4_c10_r0_io_s;
  assign ft_s5_c11_r1_io_a = fa_s4_c10_r0_io_co;
  assign fa_s6_c10_r0_io_a = ft_s5_c10_r0_io_s;
  assign fa_s6_c10_r0_io_b = ft_s5_c10_r1_io_s;
  assign ft_s7_c10_r0_io_a = fa_s6_c10_r0_io_s;
  assign ft_s7_c11_r1_io_a = fa_s6_c10_r0_io_co;
  assign ft_s8_c10_r0_io_a = ft_s7_c10_r0_io_s;
  assign io_augend[10] = ft_s8_c10_r0_io_s;
  assign fa_s1_c11_r0_io_a = fa_s0_c11_r0_io_s;
  assign fa_s1_c12_r1_io_ci = fa_s0_c11_r0_io_co;
  assign fa_s1_c11_r0_io_b = fa_s0_c11_r1_io_s;
  assign fa_s1_c12_r2_io_a = fa_s0_c11_r1_io_co;
  assign fa_s1_c11_r0_io_ci = fa_s0_c11_r2_io_s;
  assign fa_s1_c12_r2_io_b = fa_s0_c11_r2_io_co;
  assign fa_s1_c11_r1_io_a = fa_s0_c11_r3_io_s;
  assign fa_s1_c12_r2_io_ci = fa_s0_c11_r3_io_co;
  assign fa_s2_c11_r0_io_a = fa_s1_c11_r0_io_s;
  assign ft_s2_c12_r1_io_a = fa_s1_c11_r0_io_co;
  assign fa_s2_c11_r0_io_b = fa_s1_c11_r1_io_s;
  assign ft_s2_c12_r2_io_a = fa_s1_c11_r1_io_co;
  assign fa_s2_c11_r0_io_ci = ft_s1_c11_r2_io_s;
  assign fa_s3_c11_r0_io_a = fa_s2_c11_r0_io_s;
  assign ft_s3_c12_r1_io_a = fa_s2_c11_r0_io_co;
  assign fa_s3_c11_r0_io_b = ha_s2_c11_r1_io_s;
  assign ft_s3_c12_r2_io_a = ha_s2_c11_r1_io_co;
  assign ha_s4_c11_r0_io_a = fa_s3_c11_r0_io_s;
  assign ft_s4_c12_r1_io_a = fa_s3_c11_r0_io_co;
  assign ha_s4_c11_r0_io_b = ft_s3_c11_r1_io_s;
  assign ha_s5_c11_r0_io_a = ha_s4_c11_r0_io_s;
  assign fa_s5_c12_r0_io_ci = ha_s4_c11_r0_io_co;
  assign ha_s5_c11_r0_io_b = ft_s4_c11_r1_io_s;
  assign ha_s6_c11_r0_io_a = ha_s5_c11_r0_io_s;
  assign ft_s6_c12_r1_io_a = ha_s5_c11_r0_io_co;
  assign ha_s6_c11_r0_io_b = ft_s5_c11_r1_io_s;
  assign ft_s7_c11_r0_io_a = ha_s6_c11_r0_io_s;
  assign fa_s7_c12_r0_io_ci = ha_s6_c11_r0_io_co;
  assign ft_s8_c11_r0_io_a = ft_s7_c11_r0_io_s;
  assign ft_s8_c11_r1_io_a = ft_s7_c11_r1_io_s;
  assign io_augend[11] = ft_s8_c11_r0_io_s;
  assign io_addend[11] = ft_s8_c11_r1_io_s;
  assign fa_s1_c12_r0_io_a = fa_s0_c12_r0_io_s;
  assign fa_s1_c13_r2_io_a = fa_s0_c12_r0_io_co;
  assign fa_s1_c12_r0_io_b = fa_s0_c12_r1_io_s;
  assign fa_s1_c13_r2_io_b = fa_s0_c12_r1_io_co;
  assign fa_s1_c12_r0_io_ci = fa_s0_c12_r2_io_s;
  assign fa_s1_c13_r2_io_ci = fa_s0_c12_r2_io_co;
  assign fa_s1_c12_r1_io_a = fa_s0_c12_r3_io_s;
  assign ft_s1_c13_r3_io_a = fa_s0_c12_r3_io_co;
  assign fa_s1_c12_r1_io_b = ft_s0_c12_r4_io_s;
  assign fa_s2_c12_r0_io_a = fa_s1_c12_r0_io_s;
  assign fa_s2_c13_r1_io_b = fa_s1_c12_r0_io_co;
  assign fa_s2_c12_r0_io_b = fa_s1_c12_r1_io_s;
  assign fa_s2_c13_r1_io_ci = fa_s1_c12_r1_io_co;
  assign fa_s2_c12_r0_io_ci = fa_s1_c12_r2_io_s;
  assign ft_s2_c13_r2_io_a = fa_s1_c12_r2_io_co;
  assign fa_s3_c12_r0_io_a = fa_s2_c12_r0_io_s;
  assign ft_s3_c13_r1_io_a = fa_s2_c12_r0_io_co;
  assign fa_s3_c12_r0_io_b = ft_s2_c12_r1_io_s;
  assign fa_s3_c12_r0_io_ci = ft_s2_c12_r2_io_s;
  assign fa_s4_c12_r0_io_a = fa_s3_c12_r0_io_s;
  assign fa_s4_c13_r0_io_ci = fa_s3_c12_r0_io_co;
  assign fa_s4_c12_r0_io_b = ft_s3_c12_r1_io_s;
  assign fa_s4_c12_r0_io_ci = ft_s3_c12_r2_io_s;
  assign fa_s5_c12_r0_io_a = fa_s4_c12_r0_io_s;
  assign ft_s5_c13_r1_io_a = fa_s4_c12_r0_io_co;
  assign fa_s5_c12_r0_io_b = ft_s4_c12_r1_io_s;
  assign ft_s6_c12_r0_io_a = fa_s5_c12_r0_io_s;
  assign fa_s6_c13_r0_io_ci = fa_s5_c12_r0_io_co;
  assign fa_s7_c12_r0_io_a = ft_s6_c12_r0_io_s;
  assign fa_s7_c12_r0_io_b = ft_s6_c12_r1_io_s;
  assign ft_s8_c12_r0_io_a = fa_s7_c12_r0_io_s;
  assign ft_s8_c13_r1_io_a = fa_s7_c12_r0_io_co;
  assign io_augend[12] = ft_s8_c12_r0_io_s;
  assign fa_s1_c13_r0_io_a = fa_s0_c13_r0_io_s;
  assign fa_s1_c14_r1_io_ci = fa_s0_c13_r0_io_co;
  assign fa_s1_c13_r0_io_b = fa_s0_c13_r1_io_s;
  assign fa_s1_c14_r2_io_a = fa_s0_c13_r1_io_co;
  assign fa_s1_c13_r0_io_ci = fa_s0_c13_r2_io_s;
  assign fa_s1_c14_r2_io_b = fa_s0_c13_r2_io_co;
  assign fa_s1_c13_r1_io_a = fa_s0_c13_r3_io_s;
  assign fa_s1_c14_r2_io_ci = fa_s0_c13_r3_io_co;
  assign fa_s1_c13_r1_io_b = ft_s0_c13_r4_io_s;
  assign fa_s1_c13_r1_io_ci = ft_s0_c13_r5_io_s;
  assign fa_s2_c13_r0_io_a = fa_s1_c13_r0_io_s;
  assign fa_s2_c14_r1_io_a = fa_s1_c13_r0_io_co;
  assign fa_s2_c13_r0_io_b = fa_s1_c13_r1_io_s;
  assign fa_s2_c14_r1_io_b = fa_s1_c13_r1_io_co;
  assign fa_s2_c13_r0_io_ci = fa_s1_c13_r2_io_s;
  assign fa_s2_c14_r1_io_ci = fa_s1_c13_r2_io_co;
  assign fa_s2_c13_r1_io_a = ft_s1_c13_r3_io_s;
  assign fa_s3_c13_r0_io_a = fa_s2_c13_r0_io_s;
  assign fa_s3_c14_r0_io_ci = fa_s2_c13_r0_io_co;
  assign fa_s3_c13_r0_io_b = fa_s2_c13_r1_io_s;
  assign ft_s3_c14_r1_io_a = fa_s2_c13_r1_io_co;
  assign fa_s3_c13_r0_io_ci = ft_s2_c13_r2_io_s;
  assign fa_s4_c13_r0_io_a = fa_s3_c13_r0_io_s;
  assign fa_s4_c14_r0_io_ci = fa_s3_c13_r0_io_co;
  assign fa_s4_c13_r0_io_b = ft_s3_c13_r1_io_s;
  assign ft_s5_c13_r0_io_a = fa_s4_c13_r0_io_s;
  assign ft_s5_c14_r1_io_a = fa_s4_c13_r0_io_co;
  assign fa_s6_c13_r0_io_a = ft_s5_c13_r0_io_s;
  assign fa_s6_c13_r0_io_b = ft_s5_c13_r1_io_s;
  assign ft_s7_c13_r0_io_a = fa_s6_c13_r0_io_s;
  assign fa_s7_c14_r0_io_ci = fa_s6_c13_r0_io_co;
  assign ft_s8_c13_r0_io_a = ft_s7_c13_r0_io_s;
  assign io_augend[13] = ft_s8_c13_r0_io_s;
  assign io_addend[13] = ft_s8_c13_r1_io_s;
  assign fa_s1_c14_r0_io_a = fa_s0_c14_r0_io_s;
  assign fa_s1_c15_r2_io_a = fa_s0_c14_r0_io_co;
  assign fa_s1_c14_r0_io_b = fa_s0_c14_r1_io_s;
  assign fa_s1_c15_r2_io_b = fa_s0_c14_r1_io_co;
  assign fa_s1_c14_r0_io_ci = fa_s0_c14_r2_io_s;
  assign fa_s1_c15_r2_io_ci = fa_s0_c14_r2_io_co;
  assign fa_s1_c14_r1_io_a = fa_s0_c14_r3_io_s;
  assign ha_s1_c15_r3_io_a = fa_s0_c14_r3_io_co;
  assign fa_s1_c14_r1_io_b = fa_s0_c14_r4_io_s;
  assign ha_s1_c15_r3_io_b = fa_s0_c14_r4_io_co;
  assign fa_s2_c14_r0_io_a = fa_s1_c14_r0_io_s;
  assign fa_s2_c15_r1_io_b = fa_s1_c14_r0_io_co;
  assign fa_s2_c14_r0_io_b = fa_s1_c14_r1_io_s;
  assign fa_s2_c15_r1_io_ci = fa_s1_c14_r1_io_co;
  assign fa_s2_c14_r0_io_ci = fa_s1_c14_r2_io_s;
  assign ft_s2_c15_r2_io_a = fa_s1_c14_r2_io_co;
  assign fa_s3_c14_r0_io_a = fa_s2_c14_r0_io_s;
  assign ft_s3_c15_r1_io_a = fa_s2_c14_r0_io_co;
  assign fa_s3_c14_r0_io_b = fa_s2_c14_r1_io_s;
  assign ft_s3_c15_r2_io_a = fa_s2_c14_r1_io_co;
  assign fa_s4_c14_r0_io_a = fa_s3_c14_r0_io_s;
  assign ft_s4_c15_r1_io_a = fa_s3_c14_r0_io_co;
  assign fa_s4_c14_r0_io_b = ft_s3_c14_r1_io_s;
  assign ft_s5_c14_r0_io_a = fa_s4_c14_r0_io_s;
  assign fa_s5_c15_r0_io_ci = fa_s4_c14_r0_io_co;
  assign ft_s6_c14_r0_io_a = ft_s5_c14_r0_io_s;
  assign ft_s6_c14_r1_io_a = ft_s5_c14_r1_io_s;
  assign fa_s7_c14_r0_io_a = ft_s6_c14_r0_io_s;
  assign fa_s7_c14_r0_io_b = ft_s6_c14_r1_io_s;
  assign ft_s8_c14_r0_io_a = fa_s7_c14_r0_io_s;
  assign ft_s8_c15_r1_io_a = fa_s7_c14_r0_io_co;
  assign io_augend[14] = ft_s8_c14_r0_io_s;
  assign fa_s1_c15_r0_io_a = fa_s0_c15_r0_io_s;
  assign fa_s1_c16_r1_io_ci = fa_s0_c15_r0_io_co;
  assign fa_s1_c15_r0_io_b = fa_s0_c15_r1_io_s;
  assign fa_s1_c16_r2_io_a = fa_s0_c15_r1_io_co;
  assign fa_s1_c15_r0_io_ci = fa_s0_c15_r2_io_s;
  assign fa_s1_c16_r2_io_b = fa_s0_c15_r2_io_co;
  assign fa_s1_c15_r1_io_a = fa_s0_c15_r3_io_s;
  assign fa_s1_c16_r2_io_ci = fa_s0_c15_r3_io_co;
  assign fa_s1_c15_r1_io_b = fa_s0_c15_r4_io_s;
  assign ft_s1_c16_r3_io_a = fa_s0_c15_r4_io_co;
  assign fa_s1_c15_r1_io_ci = ft_s0_c15_r5_io_s;
  assign fa_s2_c15_r0_io_a = fa_s1_c15_r0_io_s;
  assign fa_s2_c16_r1_io_b = fa_s1_c15_r0_io_co;
  assign fa_s2_c15_r0_io_b = fa_s1_c15_r1_io_s;
  assign fa_s2_c16_r1_io_ci = fa_s1_c15_r1_io_co;
  assign fa_s2_c15_r0_io_ci = fa_s1_c15_r2_io_s;
  assign ha_s2_c16_r2_io_a = fa_s1_c15_r2_io_co;
  assign fa_s2_c15_r1_io_a = ha_s1_c15_r3_io_s;
  assign ha_s2_c16_r2_io_b = ha_s1_c15_r3_io_co;
  assign fa_s3_c15_r0_io_a = fa_s2_c15_r0_io_s;
  assign ft_s3_c16_r1_io_a = fa_s2_c15_r0_io_co;
  assign fa_s3_c15_r0_io_b = fa_s2_c15_r1_io_s;
  assign ft_s3_c16_r2_io_a = fa_s2_c15_r1_io_co;
  assign fa_s3_c15_r0_io_ci = ft_s2_c15_r2_io_s;
  assign fa_s4_c15_r0_io_a = fa_s3_c15_r0_io_s;
  assign ft_s4_c16_r1_io_a = fa_s3_c15_r0_io_co;
  assign fa_s4_c15_r0_io_b = ft_s3_c15_r1_io_s;
  assign fa_s4_c15_r0_io_ci = ft_s3_c15_r2_io_s;
  assign fa_s5_c15_r0_io_a = fa_s4_c15_r0_io_s;
  assign fa_s5_c16_r0_io_ci = fa_s4_c15_r0_io_co;
  assign fa_s5_c15_r0_io_b = ft_s4_c15_r1_io_s;
  assign ft_s6_c15_r0_io_a = fa_s5_c15_r0_io_s;
  assign ft_s6_c16_r1_io_a = fa_s5_c15_r0_io_co;
  assign ft_s7_c15_r0_io_a = ft_s6_c15_r0_io_s;
  assign ft_s8_c15_r0_io_a = ft_s7_c15_r0_io_s;
  assign io_augend[15] = ft_s8_c15_r0_io_s;
  assign io_addend[15] = ft_s8_c15_r1_io_s;
  assign fa_s1_c16_r0_io_a = fa_s0_c16_r0_io_s;
  assign fa_s1_c17_r2_io_a = fa_s0_c16_r0_io_co;
  assign fa_s1_c16_r0_io_b = fa_s0_c16_r1_io_s;
  assign fa_s1_c17_r2_io_b = fa_s0_c16_r1_io_co;
  assign fa_s1_c16_r0_io_ci = fa_s0_c16_r2_io_s;
  assign fa_s1_c17_r2_io_ci = fa_s0_c16_r2_io_co;
  assign fa_s1_c16_r1_io_a = fa_s0_c16_r3_io_s;
  assign ft_s1_c17_r3_io_a = fa_s0_c16_r3_io_co;
  assign fa_s1_c16_r1_io_b = fa_s0_c16_r4_io_s;
  assign ft_s1_c17_r4_io_a = fa_s0_c16_r4_io_co;
  assign fa_s2_c16_r0_io_a = fa_s1_c16_r0_io_s;
  assign fa_s2_c17_r1_io_ci = fa_s1_c16_r0_io_co;
  assign fa_s2_c16_r0_io_b = fa_s1_c16_r1_io_s;
  assign ft_s2_c17_r2_io_a = fa_s1_c16_r1_io_co;
  assign fa_s2_c16_r0_io_ci = fa_s1_c16_r2_io_s;
  assign ft_s2_c17_r3_io_a = fa_s1_c16_r2_io_co;
  assign fa_s2_c16_r1_io_a = ft_s1_c16_r3_io_s;
  assign fa_s3_c16_r0_io_a = fa_s2_c16_r0_io_s;
  assign fa_s3_c17_r1_io_b = fa_s2_c16_r0_io_co;
  assign fa_s3_c16_r0_io_b = fa_s2_c16_r1_io_s;
  assign fa_s3_c17_r1_io_ci = fa_s2_c16_r1_io_co;
  assign fa_s3_c16_r0_io_ci = ha_s2_c16_r2_io_s;
  assign ft_s3_c17_r2_io_a = ha_s2_c16_r2_io_co;
  assign fa_s4_c16_r0_io_a = fa_s3_c16_r0_io_s;
  assign ft_s4_c17_r1_io_a = fa_s3_c16_r0_io_co;
  assign fa_s4_c16_r0_io_b = ft_s3_c16_r1_io_s;
  assign fa_s4_c16_r0_io_ci = ft_s3_c16_r2_io_s;
  assign fa_s5_c16_r0_io_a = fa_s4_c16_r0_io_s;
  assign fa_s5_c17_r0_io_ci = fa_s4_c16_r0_io_co;
  assign fa_s5_c16_r0_io_b = ft_s4_c16_r1_io_s;
  assign ft_s6_c16_r0_io_a = fa_s5_c16_r0_io_s;
  assign ft_s6_c17_r1_io_a = fa_s5_c16_r0_io_co;
  assign ft_s7_c16_r0_io_a = ft_s6_c16_r0_io_s;
  assign ft_s7_c16_r1_io_a = ft_s6_c16_r1_io_s;
  assign ft_s8_c16_r0_io_a = ft_s7_c16_r0_io_s;
  assign ft_s8_c16_r1_io_a = ft_s7_c16_r1_io_s;
  assign io_augend[16] = ft_s8_c16_r0_io_s;
  assign io_addend[16] = ft_s8_c16_r1_io_s;
  assign fa_s1_c17_r0_io_a = fa_s0_c17_r0_io_s;
  assign fa_s1_c18_r1_io_ci = fa_s0_c17_r0_io_co;
  assign fa_s1_c17_r0_io_b = fa_s0_c17_r1_io_s;
  assign fa_s1_c18_r2_io_a = fa_s0_c17_r1_io_co;
  assign fa_s1_c17_r0_io_ci = fa_s0_c17_r2_io_s;
  assign fa_s1_c18_r2_io_b = fa_s0_c17_r2_io_co;
  assign fa_s1_c17_r1_io_a = fa_s0_c17_r3_io_s;
  assign fa_s1_c18_r2_io_ci = fa_s0_c17_r3_io_co;
  assign fa_s1_c17_r1_io_b = ft_s0_c17_r4_io_s;
  assign fa_s1_c17_r1_io_ci = ft_s0_c17_r5_io_s;
  assign fa_s2_c17_r0_io_a = fa_s1_c17_r0_io_s;
  assign fa_s2_c18_r1_io_a = fa_s1_c17_r0_io_co;
  assign fa_s2_c17_r0_io_b = fa_s1_c17_r1_io_s;
  assign fa_s2_c18_r1_io_b = fa_s1_c17_r1_io_co;
  assign fa_s2_c17_r0_io_ci = fa_s1_c17_r2_io_s;
  assign fa_s2_c18_r1_io_ci = fa_s1_c17_r2_io_co;
  assign fa_s2_c17_r1_io_a = ft_s1_c17_r3_io_s;
  assign fa_s2_c17_r1_io_b = ft_s1_c17_r4_io_s;
  assign fa_s3_c17_r0_io_a = fa_s2_c17_r0_io_s;
  assign fa_s3_c18_r0_io_ci = fa_s2_c17_r0_io_co;
  assign fa_s3_c17_r0_io_b = fa_s2_c17_r1_io_s;
  assign ft_s3_c18_r1_io_a = fa_s2_c17_r1_io_co;
  assign fa_s3_c17_r0_io_ci = ft_s2_c17_r2_io_s;
  assign fa_s3_c17_r1_io_a = ft_s2_c17_r3_io_s;
  assign fa_s4_c17_r0_io_a = fa_s3_c17_r0_io_s;
  assign fa_s4_c18_r0_io_ci = fa_s3_c17_r0_io_co;
  assign fa_s4_c17_r0_io_b = fa_s3_c17_r1_io_s;
  assign ft_s4_c18_r1_io_a = fa_s3_c17_r1_io_co;
  assign fa_s4_c17_r0_io_ci = ft_s3_c17_r2_io_s;
  assign fa_s5_c17_r0_io_a = fa_s4_c17_r0_io_s;
  assign fa_s5_c18_r0_io_ci = fa_s4_c17_r0_io_co;
  assign fa_s5_c17_r0_io_b = ft_s4_c17_r1_io_s;
  assign ft_s6_c17_r0_io_a = fa_s5_c17_r0_io_s;
  assign ft_s6_c18_r1_io_a = fa_s5_c17_r0_io_co;
  assign ft_s7_c17_r0_io_a = ft_s6_c17_r0_io_s;
  assign ft_s7_c17_r1_io_a = ft_s6_c17_r1_io_s;
  assign ft_s8_c17_r0_io_a = ft_s7_c17_r0_io_s;
  assign ft_s8_c17_r1_io_a = ft_s7_c17_r1_io_s;
  assign io_augend[17] = ft_s8_c17_r0_io_s;
  assign io_addend[17] = ft_s8_c17_r1_io_s;
  assign fa_s1_c18_r0_io_a = fa_s0_c18_r0_io_s;
  assign fa_s1_c19_r1_io_b = fa_s0_c18_r0_io_co;
  assign fa_s1_c18_r0_io_b = fa_s0_c18_r1_io_s;
  assign fa_s1_c19_r1_io_ci = fa_s0_c18_r1_io_co;
  assign fa_s1_c18_r0_io_ci = fa_s0_c18_r2_io_s;
  assign ha_s1_c19_r2_io_a = fa_s0_c18_r2_io_co;
  assign fa_s1_c18_r1_io_a = fa_s0_c18_r3_io_s;
  assign ha_s1_c19_r2_io_b = fa_s0_c18_r3_io_co;
  assign fa_s1_c18_r1_io_b = ft_s0_c18_r4_io_s;
  assign fa_s2_c18_r0_io_a = fa_s1_c18_r0_io_s;
  assign fa_s2_c19_r1_io_a = fa_s1_c18_r0_io_co;
  assign fa_s2_c18_r0_io_b = fa_s1_c18_r1_io_s;
  assign fa_s2_c19_r1_io_b = fa_s1_c18_r1_io_co;
  assign fa_s2_c18_r0_io_ci = fa_s1_c18_r2_io_s;
  assign fa_s2_c19_r1_io_ci = fa_s1_c18_r2_io_co;
  assign fa_s3_c18_r0_io_a = fa_s2_c18_r0_io_s;
  assign fa_s3_c19_r0_io_ci = fa_s2_c18_r0_io_co;
  assign fa_s3_c18_r0_io_b = fa_s2_c18_r1_io_s;
  assign ft_s3_c19_r1_io_a = fa_s2_c18_r1_io_co;
  assign fa_s4_c18_r0_io_a = fa_s3_c18_r0_io_s;
  assign fa_s4_c19_r0_io_ci = fa_s3_c18_r0_io_co;
  assign fa_s4_c18_r0_io_b = ft_s3_c18_r1_io_s;
  assign fa_s5_c18_r0_io_a = fa_s4_c18_r0_io_s;
  assign ft_s5_c19_r1_io_a = fa_s4_c18_r0_io_co;
  assign fa_s5_c18_r0_io_b = ft_s4_c18_r1_io_s;
  assign ft_s6_c18_r0_io_a = fa_s5_c18_r0_io_s;
  assign fa_s6_c19_r0_io_ci = fa_s5_c18_r0_io_co;
  assign ft_s7_c18_r0_io_a = ft_s6_c18_r0_io_s;
  assign ft_s7_c18_r1_io_a = ft_s6_c18_r1_io_s;
  assign ft_s8_c18_r0_io_a = ft_s7_c18_r0_io_s;
  assign ft_s8_c18_r1_io_a = ft_s7_c18_r1_io_s;
  assign io_augend[18] = ft_s8_c18_r0_io_s;
  assign io_addend[18] = ft_s8_c18_r1_io_s;
  assign fa_s1_c19_r0_io_a = fa_s0_c19_r0_io_s;
  assign fa_s1_c20_r1_io_b = fa_s0_c19_r0_io_co;
  assign fa_s1_c19_r0_io_b = fa_s0_c19_r1_io_s;
  assign fa_s1_c20_r1_io_ci = fa_s0_c19_r1_io_co;
  assign fa_s1_c19_r0_io_ci = fa_s0_c19_r2_io_s;
  assign ft_s1_c20_r2_io_a = fa_s0_c19_r2_io_co;
  assign fa_s1_c19_r1_io_a = fa_s0_c19_r3_io_s;
  assign ft_s1_c20_r3_io_a = fa_s0_c19_r3_io_co;
  assign fa_s2_c19_r0_io_a = fa_s1_c19_r0_io_s;
  assign fa_s2_c20_r1_io_b = fa_s1_c19_r0_io_co;
  assign fa_s2_c19_r0_io_b = fa_s1_c19_r1_io_s;
  assign fa_s2_c20_r1_io_ci = fa_s1_c19_r1_io_co;
  assign fa_s2_c19_r0_io_ci = ha_s1_c19_r2_io_s;
  assign ft_s2_c20_r2_io_a = ha_s1_c19_r2_io_co;
  assign fa_s3_c19_r0_io_a = fa_s2_c19_r0_io_s;
  assign ft_s3_c20_r1_io_a = fa_s2_c19_r0_io_co;
  assign fa_s3_c19_r0_io_b = fa_s2_c19_r1_io_s;
  assign ft_s3_c20_r2_io_a = fa_s2_c19_r1_io_co;
  assign fa_s4_c19_r0_io_a = fa_s3_c19_r0_io_s;
  assign ft_s4_c20_r1_io_a = fa_s3_c19_r0_io_co;
  assign fa_s4_c19_r0_io_b = ft_s3_c19_r1_io_s;
  assign ft_s5_c19_r0_io_a = fa_s4_c19_r0_io_s;
  assign fa_s5_c20_r0_io_ci = fa_s4_c19_r0_io_co;
  assign fa_s6_c19_r0_io_a = ft_s5_c19_r0_io_s;
  assign fa_s6_c19_r0_io_b = ft_s5_c19_r1_io_s;
  assign ft_s7_c19_r0_io_a = fa_s6_c19_r0_io_s;
  assign ft_s7_c20_r1_io_a = fa_s6_c19_r0_io_co;
  assign ft_s8_c19_r0_io_a = ft_s7_c19_r0_io_s;
  assign io_augend[19] = ft_s8_c19_r0_io_s;
  assign fa_s1_c20_r0_io_a = fa_s0_c20_r0_io_s;
  assign fa_s1_c21_r1_io_b = fa_s0_c20_r0_io_co;
  assign fa_s1_c20_r0_io_b = fa_s0_c20_r1_io_s;
  assign fa_s1_c21_r1_io_ci = fa_s0_c20_r1_io_co;
  assign fa_s1_c20_r0_io_ci = fa_s0_c20_r2_io_s;
  assign ha_s1_c21_r2_io_a = fa_s0_c20_r2_io_co;
  assign fa_s1_c20_r1_io_a = ha_s0_c20_r3_io_s;
  assign ha_s1_c21_r2_io_b = ha_s0_c20_r3_io_co;
  assign fa_s2_c20_r0_io_a = fa_s1_c20_r0_io_s;
  assign ft_s2_c21_r1_io_a = fa_s1_c20_r0_io_co;
  assign fa_s2_c20_r0_io_b = fa_s1_c20_r1_io_s;
  assign ft_s2_c21_r2_io_a = fa_s1_c20_r1_io_co;
  assign fa_s2_c20_r0_io_ci = ft_s1_c20_r2_io_s;
  assign fa_s2_c20_r1_io_a = ft_s1_c20_r3_io_s;
  assign fa_s3_c20_r0_io_a = fa_s2_c20_r0_io_s;
  assign ft_s3_c21_r1_io_a = fa_s2_c20_r0_io_co;
  assign fa_s3_c20_r0_io_b = fa_s2_c20_r1_io_s;
  assign ft_s3_c21_r2_io_a = fa_s2_c20_r1_io_co;
  assign fa_s3_c20_r0_io_ci = ft_s2_c20_r2_io_s;
  assign fa_s4_c20_r0_io_a = fa_s3_c20_r0_io_s;
  assign ft_s4_c21_r1_io_a = fa_s3_c20_r0_io_co;
  assign fa_s4_c20_r0_io_b = ft_s3_c20_r1_io_s;
  assign fa_s4_c20_r0_io_ci = ft_s3_c20_r2_io_s;
  assign fa_s5_c20_r0_io_a = fa_s4_c20_r0_io_s;
  assign fa_s5_c21_r0_io_ci = fa_s4_c20_r0_io_co;
  assign fa_s5_c20_r0_io_b = ft_s4_c20_r1_io_s;
  assign ft_s6_c20_r0_io_a = fa_s5_c20_r0_io_s;
  assign ft_s6_c21_r1_io_a = fa_s5_c20_r0_io_co;
  assign ft_s7_c20_r0_io_a = ft_s6_c20_r0_io_s;
  assign ft_s8_c20_r0_io_a = ft_s7_c20_r0_io_s;
  assign ft_s8_c20_r1_io_a = ft_s7_c20_r1_io_s;
  assign io_augend[20] = ft_s8_c20_r0_io_s;
  assign io_addend[20] = ft_s8_c20_r1_io_s;
  assign fa_s1_c21_r0_io_a = fa_s0_c21_r0_io_s;
  assign fa_s1_c22_r1_io_a = fa_s0_c21_r0_io_co;
  assign fa_s1_c21_r0_io_b = fa_s0_c21_r1_io_s;
  assign fa_s1_c22_r1_io_b = fa_s0_c21_r1_io_co;
  assign fa_s1_c21_r0_io_ci = fa_s0_c21_r2_io_s;
  assign fa_s1_c22_r1_io_ci = fa_s0_c21_r2_io_co;
  assign fa_s1_c21_r1_io_a = ft_s0_c21_r3_io_s;
  assign fa_s2_c21_r0_io_a = fa_s1_c21_r0_io_s;
  assign fa_s2_c22_r0_io_ci = fa_s1_c21_r0_io_co;
  assign fa_s2_c21_r0_io_b = fa_s1_c21_r1_io_s;
  assign ha_s2_c22_r1_io_a = fa_s1_c21_r1_io_co;
  assign fa_s2_c21_r0_io_ci = ha_s1_c21_r2_io_s;
  assign ha_s2_c22_r1_io_b = ha_s1_c21_r2_io_co;
  assign fa_s3_c21_r0_io_a = fa_s2_c21_r0_io_s;
  assign fa_s3_c22_r0_io_ci = fa_s2_c21_r0_io_co;
  assign fa_s3_c21_r0_io_b = ft_s2_c21_r1_io_s;
  assign fa_s3_c21_r0_io_ci = ft_s2_c21_r2_io_s;
  assign fa_s4_c21_r0_io_a = fa_s3_c21_r0_io_s;
  assign ft_s4_c22_r1_io_a = fa_s3_c21_r0_io_co;
  assign fa_s4_c21_r0_io_b = ft_s3_c21_r1_io_s;
  assign fa_s4_c21_r0_io_ci = ft_s3_c21_r2_io_s;
  assign fa_s5_c21_r0_io_a = fa_s4_c21_r0_io_s;
  assign fa_s5_c22_r0_io_ci = fa_s4_c21_r0_io_co;
  assign fa_s5_c21_r0_io_b = ft_s4_c21_r1_io_s;
  assign ft_s6_c21_r0_io_a = fa_s5_c21_r0_io_s;
  assign ft_s6_c22_r1_io_a = fa_s5_c21_r0_io_co;
  assign ft_s7_c21_r0_io_a = ft_s6_c21_r0_io_s;
  assign ft_s7_c21_r1_io_a = ft_s6_c21_r1_io_s;
  assign ft_s8_c21_r0_io_a = ft_s7_c21_r0_io_s;
  assign ft_s8_c21_r1_io_a = ft_s7_c21_r1_io_s;
  assign io_augend[21] = ft_s8_c21_r0_io_s;
  assign io_addend[21] = ft_s8_c21_r1_io_s;
  assign fa_s1_c22_r0_io_a = fa_s0_c22_r0_io_s;
  assign fa_s1_c23_r1_io_b = fa_s0_c22_r0_io_co;
  assign fa_s1_c22_r0_io_b = fa_s0_c22_r1_io_s;
  assign fa_s1_c23_r1_io_ci = fa_s0_c22_r1_io_co;
  assign fa_s1_c22_r0_io_ci = fa_s0_c22_r2_io_s;
  assign ft_s1_c23_r2_io_a = fa_s0_c22_r2_io_co;
  assign fa_s2_c22_r0_io_a = fa_s1_c22_r0_io_s;
  assign ft_s2_c23_r1_io_a = fa_s1_c22_r0_io_co;
  assign fa_s2_c22_r0_io_b = fa_s1_c22_r1_io_s;
  assign ft_s2_c23_r2_io_a = fa_s1_c22_r1_io_co;
  assign fa_s3_c22_r0_io_a = fa_s2_c22_r0_io_s;
  assign ft_s3_c23_r1_io_a = fa_s2_c22_r0_io_co;
  assign fa_s3_c22_r0_io_b = ha_s2_c22_r1_io_s;
  assign ft_s3_c23_r2_io_a = ha_s2_c22_r1_io_co;
  assign ft_s4_c22_r0_io_a = fa_s3_c22_r0_io_s;
  assign ft_s4_c23_r1_io_a = fa_s3_c22_r0_io_co;
  assign fa_s5_c22_r0_io_a = ft_s4_c22_r0_io_s;
  assign fa_s5_c22_r0_io_b = ft_s4_c22_r1_io_s;
  assign ft_s6_c22_r0_io_a = fa_s5_c22_r0_io_s;
  assign fa_s6_c23_r0_io_ci = fa_s5_c22_r0_io_co;
  assign ft_s7_c22_r0_io_a = ft_s6_c22_r0_io_s;
  assign ft_s7_c22_r1_io_a = ft_s6_c22_r1_io_s;
  assign ft_s8_c22_r0_io_a = ft_s7_c22_r0_io_s;
  assign ft_s8_c22_r1_io_a = ft_s7_c22_r1_io_s;
  assign io_augend[22] = ft_s8_c22_r0_io_s;
  assign io_addend[22] = ft_s8_c22_r1_io_s;
  assign fa_s1_c23_r0_io_a = fa_s0_c23_r0_io_s;
  assign ft_s1_c24_r1_io_a = fa_s0_c23_r0_io_co;
  assign fa_s1_c23_r0_io_b = fa_s0_c23_r1_io_s;
  assign ft_s1_c24_r2_io_a = fa_s0_c23_r1_io_co;
  assign fa_s1_c23_r0_io_ci = ft_s0_c23_r2_io_s;
  assign fa_s1_c23_r1_io_a = ft_s0_c23_r3_io_s;
  assign fa_s2_c23_r0_io_a = fa_s1_c23_r0_io_s;
  assign ft_s2_c24_r1_io_a = fa_s1_c23_r0_io_co;
  assign fa_s2_c23_r0_io_b = fa_s1_c23_r1_io_s;
  assign ft_s2_c24_r2_io_a = fa_s1_c23_r1_io_co;
  assign fa_s2_c23_r0_io_ci = ft_s1_c23_r2_io_s;
  assign fa_s3_c23_r0_io_a = fa_s2_c23_r0_io_s;
  assign ft_s3_c24_r1_io_a = fa_s2_c23_r0_io_co;
  assign fa_s3_c23_r0_io_b = ft_s2_c23_r1_io_s;
  assign fa_s3_c23_r0_io_ci = ft_s2_c23_r2_io_s;
  assign fa_s4_c23_r0_io_a = fa_s3_c23_r0_io_s;
  assign fa_s4_c24_r0_io_ci = fa_s3_c23_r0_io_co;
  assign fa_s4_c23_r0_io_b = ft_s3_c23_r1_io_s;
  assign fa_s4_c23_r0_io_ci = ft_s3_c23_r2_io_s;
  assign ft_s5_c23_r0_io_a = fa_s4_c23_r0_io_s;
  assign ft_s5_c24_r1_io_a = fa_s4_c23_r0_io_co;
  assign ft_s5_c23_r1_io_a = ft_s4_c23_r1_io_s;
  assign fa_s6_c23_r0_io_a = ft_s5_c23_r0_io_s;
  assign fa_s6_c23_r0_io_b = ft_s5_c23_r1_io_s;
  assign ft_s7_c23_r0_io_a = fa_s6_c23_r0_io_s;
  assign fa_s7_c24_r0_io_ci = fa_s6_c23_r0_io_co;
  assign ft_s8_c23_r0_io_a = ft_s7_c23_r0_io_s;
  assign io_augend[23] = ft_s8_c23_r0_io_s;
  assign fa_s1_c24_r0_io_a = fa_s0_c24_r0_io_s;
  assign fa_s1_c25_r0_io_ci = fa_s0_c24_r0_io_co;
  assign fa_s1_c24_r0_io_b = fa_s0_c24_r1_io_s;
  assign ft_s1_c25_r1_io_a = fa_s0_c24_r1_io_co;
  assign fa_s1_c24_r0_io_ci = ft_s0_c24_r2_io_s;
  assign fa_s2_c24_r0_io_a = fa_s1_c24_r0_io_s;
  assign fa_s2_c25_r0_io_ci = fa_s1_c24_r0_io_co;
  assign fa_s2_c24_r0_io_b = ft_s1_c24_r1_io_s;
  assign fa_s2_c24_r0_io_ci = ft_s1_c24_r2_io_s;
  assign fa_s3_c24_r0_io_a = fa_s2_c24_r0_io_s;
  assign ha_s3_c25_r0_io_b = fa_s2_c24_r0_io_co;
  assign fa_s3_c24_r0_io_b = ft_s2_c24_r1_io_s;
  assign fa_s3_c24_r0_io_ci = ft_s2_c24_r2_io_s;
  assign fa_s4_c24_r0_io_a = fa_s3_c24_r0_io_s;
  assign ha_s4_c25_r0_io_b = fa_s3_c24_r0_io_co;
  assign fa_s4_c24_r0_io_b = ft_s3_c24_r1_io_s;
  assign ft_s5_c24_r0_io_a = fa_s4_c24_r0_io_s;
  assign ft_s5_c25_r1_io_a = fa_s4_c24_r0_io_co;
  assign ft_s6_c24_r0_io_a = ft_s5_c24_r0_io_s;
  assign ft_s6_c24_r1_io_a = ft_s5_c24_r1_io_s;
  assign fa_s7_c24_r0_io_a = ft_s6_c24_r0_io_s;
  assign fa_s7_c24_r0_io_b = ft_s6_c24_r1_io_s;
  assign ft_s8_c24_r0_io_a = fa_s7_c24_r0_io_s;
  assign fa_s8_c25_r0_io_ci = fa_s7_c24_r0_io_co;
  assign io_augend[24] = ft_s8_c24_r0_io_s;
  assign fa_s1_c25_r0_io_a = fa_s0_c25_r0_io_s;
  assign ft_s1_c26_r1_io_a = fa_s0_c25_r0_io_co;
  assign fa_s1_c25_r0_io_b = fa_s0_c25_r1_io_s;
  assign ft_s1_c26_r2_io_a = fa_s0_c25_r1_io_co;
  assign fa_s2_c25_r0_io_a = fa_s1_c25_r0_io_s;
  assign ft_s2_c26_r1_io_a = fa_s1_c25_r0_io_co;
  assign fa_s2_c25_r0_io_b = ft_s1_c25_r1_io_s;
  assign ha_s3_c25_r0_io_a = fa_s2_c25_r0_io_s;
  assign fa_s3_c26_r0_io_ci = fa_s2_c25_r0_io_co;
  assign ha_s4_c25_r0_io_a = ha_s3_c25_r0_io_s;
  assign ft_s4_c26_r1_io_a = ha_s3_c25_r0_io_co;
  assign ft_s5_c25_r0_io_a = ha_s4_c25_r0_io_s;
  assign fa_s5_c26_r0_io_ci = ha_s4_c25_r0_io_co;
  assign ft_s6_c25_r0_io_a = ft_s5_c25_r0_io_s;
  assign ft_s6_c25_r1_io_a = ft_s5_c25_r1_io_s;
  assign ft_s7_c25_r0_io_a = ft_s6_c25_r0_io_s;
  assign ft_s7_c25_r1_io_a = ft_s6_c25_r1_io_s;
  assign fa_s8_c25_r0_io_a = ft_s7_c25_r0_io_s;
  assign fa_s8_c25_r0_io_b = ft_s7_c25_r1_io_s;
  assign io_augend[25] = fa_s8_c25_r0_io_s;
  assign io_addend[26] = fa_s8_c25_r0_io_co;
  assign fa_s1_c26_r0_io_a = fa_s0_c26_r0_io_s;
  assign fa_s1_c27_r0_io_ci = fa_s0_c26_r0_io_co;
  assign fa_s1_c26_r0_io_b = ft_s0_c26_r1_io_s;
  assign fa_s1_c26_r0_io_ci = ft_s0_c26_r2_io_s;
  assign fa_s2_c26_r0_io_a = fa_s1_c26_r0_io_s;
  assign ft_s2_c27_r1_io_a = fa_s1_c26_r0_io_co;
  assign fa_s2_c26_r0_io_b = ft_s1_c26_r1_io_s;
  assign fa_s2_c26_r0_io_ci = ft_s1_c26_r2_io_s;
  assign fa_s3_c26_r0_io_a = fa_s2_c26_r0_io_s;
  assign fa_s3_c27_r0_io_ci = fa_s2_c26_r0_io_co;
  assign fa_s3_c26_r0_io_b = ft_s2_c26_r1_io_s;
  assign ft_s4_c26_r0_io_a = fa_s3_c26_r0_io_s;
  assign ft_s4_c27_r1_io_a = fa_s3_c26_r0_io_co;
  assign fa_s5_c26_r0_io_a = ft_s4_c26_r0_io_s;
  assign fa_s5_c26_r0_io_b = ft_s4_c26_r1_io_s;
  assign ft_s6_c26_r0_io_a = fa_s5_c26_r0_io_s;
  assign fa_s6_c27_r0_io_ci = fa_s5_c26_r0_io_co;
  assign ft_s7_c26_r0_io_a = ft_s6_c26_r0_io_s;
  assign ft_s8_c26_r0_io_a = ft_s7_c26_r0_io_s;
  assign io_augend[26] = ft_s8_c26_r0_io_s;
  assign fa_s1_c27_r0_io_a = fa_s0_c27_r0_io_s;
  assign ha_s1_c28_r0_io_b = fa_s0_c27_r0_io_co;
  assign fa_s1_c27_r0_io_b = ft_s0_c27_r1_io_s;
  assign ft_s2_c27_r0_io_a = fa_s1_c27_r0_io_s;
  assign ha_s2_c28_r0_io_b = fa_s1_c27_r0_io_co;
  assign fa_s3_c27_r0_io_a = ft_s2_c27_r0_io_s;
  assign fa_s3_c27_r0_io_b = ft_s2_c27_r1_io_s;
  assign ft_s4_c27_r0_io_a = fa_s3_c27_r0_io_s;
  assign ft_s4_c28_r1_io_a = fa_s3_c27_r0_io_co;
  assign ft_s5_c27_r0_io_a = ft_s4_c27_r0_io_s;
  assign ft_s5_c27_r1_io_a = ft_s4_c27_r1_io_s;
  assign fa_s6_c27_r0_io_a = ft_s5_c27_r0_io_s;
  assign fa_s6_c27_r0_io_b = ft_s5_c27_r1_io_s;
  assign ft_s7_c27_r0_io_a = fa_s6_c27_r0_io_s;
  assign fa_s7_c28_r0_io_ci = fa_s6_c27_r0_io_co;
  assign ft_s8_c27_r0_io_a = ft_s7_c27_r0_io_s;
  assign io_augend[27] = ft_s8_c27_r0_io_s;
  assign ha_s1_c28_r0_io_a = fa_s0_c28_r0_io_s;
  assign ft_s1_c29_r1_io_a = fa_s0_c28_r0_io_co;
  assign ha_s2_c28_r0_io_a = ha_s1_c28_r0_io_s;
  assign fa_s2_c29_r0_io_ci = ha_s1_c28_r0_io_co;
  assign ft_s3_c28_r0_io_a = ha_s2_c28_r0_io_s;
  assign ft_s3_c29_r1_io_a = ha_s2_c28_r0_io_co;
  assign ft_s4_c28_r0_io_a = ft_s3_c28_r0_io_s;
  assign ft_s5_c28_r0_io_a = ft_s4_c28_r0_io_s;
  assign ft_s5_c28_r1_io_a = ft_s4_c28_r1_io_s;
  assign ft_s6_c28_r0_io_a = ft_s5_c28_r0_io_s;
  assign ft_s6_c28_r1_io_a = ft_s5_c28_r1_io_s;
  assign fa_s7_c28_r0_io_a = ft_s6_c28_r0_io_s;
  assign fa_s7_c28_r0_io_b = ft_s6_c28_r1_io_s;
  assign ft_s8_c28_r0_io_a = fa_s7_c28_r0_io_s;
  assign fa_s8_c29_r0_io_ci = fa_s7_c28_r0_io_co;
  assign io_augend[28] = ft_s8_c28_r0_io_s;
  assign ft_s1_c29_r0_io_a = ha_s0_c29_r0_io_s;
  assign ft_s1_c30_r1_io_a = ha_s0_c29_r0_io_co;
  assign fa_s2_c29_r0_io_a = ft_s1_c29_r0_io_s;
  assign fa_s2_c29_r0_io_b = ft_s1_c29_r1_io_s;
  assign ft_s3_c29_r0_io_a = fa_s2_c29_r0_io_s;
  assign fa_s3_c30_r0_io_ci = fa_s2_c29_r0_io_co;
  assign ft_s4_c29_r0_io_a = ft_s3_c29_r0_io_s;
  assign ft_s4_c29_r1_io_a = ft_s3_c29_r1_io_s;
  assign ft_s5_c29_r0_io_a = ft_s4_c29_r0_io_s;
  assign ft_s5_c29_r1_io_a = ft_s4_c29_r1_io_s;
  assign ft_s6_c29_r0_io_a = ft_s5_c29_r0_io_s;
  assign ft_s6_c29_r1_io_a = ft_s5_c29_r1_io_s;
  assign ft_s7_c29_r0_io_a = ft_s6_c29_r0_io_s;
  assign ft_s7_c29_r1_io_a = ft_s6_c29_r1_io_s;
  assign fa_s8_c29_r0_io_a = ft_s7_c29_r0_io_s;
  assign fa_s8_c29_r0_io_b = ft_s7_c29_r1_io_s;
  assign io_augend[29] = fa_s8_c29_r0_io_s;
  assign io_addend[30] = fa_s8_c29_r0_io_co;
  assign ft_s1_c30_r0_io_a = ft_s0_c30_r0_io_s;
  assign ft_s2_c30_r0_io_a = ft_s1_c30_r0_io_s;
  assign ft_s2_c30_r1_io_a = ft_s1_c30_r1_io_s;
  assign fa_s3_c30_r0_io_a = ft_s2_c30_r0_io_s;
  assign fa_s3_c30_r0_io_b = ft_s2_c30_r1_io_s;
  assign ft_s4_c30_r0_io_a = fa_s3_c30_r0_io_s;
  assign ft_s4_c31_r0_io_a = fa_s3_c30_r0_io_co;
  assign ft_s5_c30_r0_io_a = ft_s4_c30_r0_io_s;
  assign ft_s6_c30_r0_io_a = ft_s5_c30_r0_io_s;
  assign ft_s7_c30_r0_io_a = ft_s6_c30_r0_io_s;
  assign ft_s8_c30_r0_io_a = ft_s7_c30_r0_io_s;
  assign io_augend[30] = ft_s8_c30_r0_io_s;
  assign ft_s5_c31_r0_io_a = ft_s4_c31_r0_io_s;
  assign ft_s6_c31_r0_io_a = ft_s5_c31_r0_io_s;
  assign ft_s7_c31_r0_io_a = ft_s6_c31_r0_io_s;
  assign ft_s8_c31_r0_io_a = ft_s7_c31_r0_io_s;
  assign io_augend[31] = ft_s8_c31_r0_io_s;
  assign io_addend[0] = 1'b0;
  assign io_addend[1] = 1'b0;
  assign io_addend[3] = 1'b0;
  assign io_addend[5] = 1'b0;
  assign io_addend[7] = 1'b0;
  assign io_addend[9] = 1'b0;
  assign io_addend[10] = 1'b0;
  assign io_addend[12] = 1'b0;
  assign io_addend[14] = 1'b0;
  assign io_addend[19] = 1'b0;
  assign io_addend[23] = 1'b0;
  assign io_addend[24] = 1'b0;
  assign io_addend[25] = 1'b0;
  assign io_addend[27] = 1'b0;
  assign io_addend[28] = 1'b0;
  assign io_addend[29] = 1'b0;
  assign io_addend[31] = 1'b0;
endmodule

`ifndef OP_PPADDER
`define OP_PPADDER

module PG(
  input   io_i_a,
  input   io_i_b,
  output  io_o_p,
  output  io_o_g
);
  assign io_o_p = io_i_a ^ io_i_b;
  assign io_o_g = io_i_a & io_i_b;
endmodule

module Black(
  input   io_i_pj,
  input   io_i_gj,
  input   io_i_pk,
  input   io_i_gk,
  output  io_o_g,
  output  io_o_p
);
  wire  _T = io_i_gj & io_i_pk;
  assign io_o_g = io_i_gk | _T;
  assign io_o_p = io_i_pk & io_i_pj;
endmodule

`endif

module CarryPropagateAdder (
  input        clock,
  input        reset,
  input  [31:0] io_augend,
  input  [31:0] io_addend,
  output [31:0] io_outs
);

  wire  PG_0_io_i_a;
  wire  PG_0_io_i_b;
  wire  PG_0_io_o_p;
  wire  PG_0_io_o_g;
  PG PG_0 (
    .io_i_a(PG_0_io_i_a),
    .io_i_b(PG_0_io_i_b),
    .io_o_p(PG_0_io_o_p),
    .io_o_g(PG_0_io_o_g)
  );

  wire  Black_1_io_i_pj;
  wire  Black_1_io_i_gj;
  wire  Black_1_io_i_pk;
  wire  Black_1_io_i_gk;
  wire  Black_1_io_o_g;
  wire  Black_1_io_o_p;
  Black Black_1 (
    .io_i_pj(Black_1_io_i_pj),
    .io_i_gj(Black_1_io_i_gj),
    .io_i_pk(Black_1_io_i_pk),
    .io_i_gk(Black_1_io_i_gk),
    .io_o_g(Black_1_io_o_g),
    .io_o_p(Black_1_io_o_p)
  );

  wire  Black_3_io_i_pj;
  wire  Black_3_io_i_gj;
  wire  Black_3_io_i_pk;
  wire  Black_3_io_i_gk;
  wire  Black_3_io_o_g;
  wire  Black_3_io_o_p;
  Black Black_3 (
    .io_i_pj(Black_3_io_i_pj),
    .io_i_gj(Black_3_io_i_gj),
    .io_i_pk(Black_3_io_i_pk),
    .io_i_gk(Black_3_io_i_gk),
    .io_o_g(Black_3_io_o_g),
    .io_o_p(Black_3_io_o_p)
  );

  wire  Black_7_io_i_pj;
  wire  Black_7_io_i_gj;
  wire  Black_7_io_i_pk;
  wire  Black_7_io_i_gk;
  wire  Black_7_io_o_g;
  wire  Black_7_io_o_p;
  Black Black_7 (
    .io_i_pj(Black_7_io_i_pj),
    .io_i_gj(Black_7_io_i_gj),
    .io_i_pk(Black_7_io_i_pk),
    .io_i_gk(Black_7_io_i_gk),
    .io_o_g(Black_7_io_o_g),
    .io_o_p(Black_7_io_o_p)
  );

  wire  Black_15_io_i_pj;
  wire  Black_15_io_i_gj;
  wire  Black_15_io_i_pk;
  wire  Black_15_io_i_gk;
  wire  Black_15_io_o_g;
  wire  Black_15_io_o_p;
  Black Black_15 (
    .io_i_pj(Black_15_io_i_pj),
    .io_i_gj(Black_15_io_i_gj),
    .io_i_pk(Black_15_io_i_pk),
    .io_i_gk(Black_15_io_i_gk),
    .io_o_g(Black_15_io_o_g),
    .io_o_p(Black_15_io_o_p)
  );

  wire  Black_31_io_i_pj;
  wire  Black_31_io_i_gj;
  wire  Black_31_io_i_pk;
  wire  Black_31_io_i_gk;
  wire  Black_31_io_o_g;
  wire  Black_31_io_o_p;
  Black Black_31 (
    .io_i_pj(Black_31_io_i_pj),
    .io_i_gj(Black_31_io_i_gj),
    .io_i_pk(Black_31_io_i_pk),
    .io_i_gk(Black_31_io_i_gk),
    .io_o_g(Black_31_io_o_g),
    .io_o_p(Black_31_io_o_p)
  );

  wire  PG_32_io_i_a;
  wire  PG_32_io_i_b;
  wire  PG_32_io_o_p;
  wire  PG_32_io_o_g;
  PG PG_32 (
    .io_i_a(PG_32_io_i_a),
    .io_i_b(PG_32_io_i_b),
    .io_o_p(PG_32_io_o_p),
    .io_o_g(PG_32_io_o_g)
  );

  wire  Black_34_io_i_pj;
  wire  Black_34_io_i_gj;
  wire  Black_34_io_i_pk;
  wire  Black_34_io_i_gk;
  wire  Black_34_io_o_g;
  wire  Black_34_io_o_p;
  Black Black_34 (
    .io_i_pj(Black_34_io_i_pj),
    .io_i_gj(Black_34_io_i_gj),
    .io_i_pk(Black_34_io_i_pk),
    .io_i_gk(Black_34_io_i_gk),
    .io_o_g(Black_34_io_o_g),
    .io_o_p(Black_34_io_o_p)
  );

  wire  Black_38_io_i_pj;
  wire  Black_38_io_i_gj;
  wire  Black_38_io_i_pk;
  wire  Black_38_io_i_gk;
  wire  Black_38_io_o_g;
  wire  Black_38_io_o_p;
  Black Black_38 (
    .io_i_pj(Black_38_io_i_pj),
    .io_i_gj(Black_38_io_i_gj),
    .io_i_pk(Black_38_io_i_pk),
    .io_i_gk(Black_38_io_i_gk),
    .io_o_g(Black_38_io_o_g),
    .io_o_p(Black_38_io_o_p)
  );

  wire  Black_46_io_i_pj;
  wire  Black_46_io_i_gj;
  wire  Black_46_io_i_pk;
  wire  Black_46_io_i_gk;
  wire  Black_46_io_o_g;
  wire  Black_46_io_o_p;
  Black Black_46 (
    .io_i_pj(Black_46_io_i_pj),
    .io_i_gj(Black_46_io_i_gj),
    .io_i_pk(Black_46_io_i_pk),
    .io_i_gk(Black_46_io_i_gk),
    .io_o_g(Black_46_io_o_g),
    .io_o_p(Black_46_io_o_p)
  );

  wire  Black_53_io_i_pj;
  wire  Black_53_io_i_gj;
  wire  Black_53_io_i_pk;
  wire  Black_53_io_i_gk;
  wire  Black_53_io_o_g;
  wire  Black_53_io_o_p;
  Black Black_53 (
    .io_i_pj(Black_53_io_i_pj),
    .io_i_gj(Black_53_io_i_gj),
    .io_i_pk(Black_53_io_i_pk),
    .io_i_gk(Black_53_io_i_gk),
    .io_o_g(Black_53_io_o_g),
    .io_o_p(Black_53_io_o_p)
  );

  wire  Black_62_io_i_pj;
  wire  Black_62_io_i_gj;
  wire  Black_62_io_i_pk;
  wire  Black_62_io_i_gk;
  wire  Black_62_io_o_g;
  wire  Black_62_io_o_p;
  Black Black_62 (
    .io_i_pj(Black_62_io_i_pj),
    .io_i_gj(Black_62_io_i_gj),
    .io_i_pk(Black_62_io_i_pk),
    .io_i_gk(Black_62_io_i_gk),
    .io_o_g(Black_62_io_o_g),
    .io_o_p(Black_62_io_o_p)
  );

  wire  PG_63_io_i_a;
  wire  PG_63_io_i_b;
  wire  PG_63_io_o_p;
  wire  PG_63_io_o_g;
  PG PG_63 (
    .io_i_a(PG_63_io_i_a),
    .io_i_b(PG_63_io_i_b),
    .io_o_p(PG_63_io_o_p),
    .io_o_g(PG_63_io_o_g)
  );

  wire  Black_64_io_i_pj;
  wire  Black_64_io_i_gj;
  wire  Black_64_io_i_pk;
  wire  Black_64_io_i_gk;
  wire  Black_64_io_o_g;
  wire  Black_64_io_o_p;
  Black Black_64 (
    .io_i_pj(Black_64_io_i_pj),
    .io_i_gj(Black_64_io_i_gj),
    .io_i_pk(Black_64_io_i_pk),
    .io_i_gk(Black_64_io_i_gk),
    .io_o_g(Black_64_io_o_g),
    .io_o_p(Black_64_io_o_p)
  );

  wire  Black_68_io_i_pj;
  wire  Black_68_io_i_gj;
  wire  Black_68_io_i_pk;
  wire  Black_68_io_i_gk;
  wire  Black_68_io_o_g;
  wire  Black_68_io_o_p;
  Black Black_68 (
    .io_i_pj(Black_68_io_i_pj),
    .io_i_gj(Black_68_io_i_gj),
    .io_i_pk(Black_68_io_i_pk),
    .io_i_gk(Black_68_io_i_gk),
    .io_o_g(Black_68_io_o_g),
    .io_o_p(Black_68_io_o_p)
  );

  wire  Black_87_io_i_pj;
  wire  Black_87_io_i_gj;
  wire  Black_87_io_i_pk;
  wire  Black_87_io_i_gk;
  wire  Black_87_io_o_g;
  wire  Black_87_io_o_p;
  Black Black_87 (
    .io_i_pj(Black_87_io_i_pj),
    .io_i_gj(Black_87_io_i_gj),
    .io_i_pk(Black_87_io_i_pk),
    .io_i_gk(Black_87_io_i_gk),
    .io_o_g(Black_87_io_o_g),
    .io_o_p(Black_87_io_o_p)
  );

  wire  Black_90_io_i_pj;
  wire  Black_90_io_i_gj;
  wire  Black_90_io_i_pk;
  wire  Black_90_io_i_gk;
  wire  Black_90_io_o_g;
  wire  Black_90_io_o_p;
  Black Black_90 (
    .io_i_pj(Black_90_io_i_pj),
    .io_i_gj(Black_90_io_i_gj),
    .io_i_pk(Black_90_io_i_pk),
    .io_i_gk(Black_90_io_i_gk),
    .io_o_g(Black_90_io_o_g),
    .io_o_p(Black_90_io_o_p)
  );

  wire  Black_92_io_i_pj;
  wire  Black_92_io_i_gj;
  wire  Black_92_io_i_pk;
  wire  Black_92_io_i_gk;
  wire  Black_92_io_o_g;
  wire  Black_92_io_o_p;
  Black Black_92 (
    .io_i_pj(Black_92_io_i_pj),
    .io_i_gj(Black_92_io_i_gj),
    .io_i_pk(Black_92_io_i_pk),
    .io_i_gk(Black_92_io_i_gk),
    .io_o_g(Black_92_io_o_g),
    .io_o_p(Black_92_io_o_p)
  );

  wire  PG_93_io_i_a;
  wire  PG_93_io_i_b;
  wire  PG_93_io_o_p;
  wire  PG_93_io_o_g;
  PG PG_93 (
    .io_i_a(PG_93_io_i_a),
    .io_i_b(PG_93_io_i_b),
    .io_o_p(PG_93_io_o_p),
    .io_o_g(PG_93_io_o_g)
  );

  wire  Black_99_io_i_pj;
  wire  Black_99_io_i_gj;
  wire  Black_99_io_i_pk;
  wire  Black_99_io_i_gk;
  wire  Black_99_io_o_g;
  wire  Black_99_io_o_p;
  Black Black_99 (
    .io_i_pj(Black_99_io_i_pj),
    .io_i_gj(Black_99_io_i_gj),
    .io_i_pk(Black_99_io_i_pk),
    .io_i_gk(Black_99_io_i_gk),
    .io_o_g(Black_99_io_o_g),
    .io_o_p(Black_99_io_o_p)
  );

  wire  Black_105_io_i_pj;
  wire  Black_105_io_i_gj;
  wire  Black_105_io_i_pk;
  wire  Black_105_io_i_gk;
  wire  Black_105_io_o_g;
  wire  Black_105_io_o_p;
  Black Black_105 (
    .io_i_pj(Black_105_io_i_pj),
    .io_i_gj(Black_105_io_i_gj),
    .io_i_pk(Black_105_io_i_pk),
    .io_i_gk(Black_105_io_i_gk),
    .io_o_g(Black_105_io_o_g),
    .io_o_p(Black_105_io_o_p)
  );

  wire  Black_121_io_i_pj;
  wire  Black_121_io_i_gj;
  wire  Black_121_io_i_pk;
  wire  Black_121_io_i_gk;
  wire  Black_121_io_o_g;
  wire  Black_121_io_o_p;
  Black Black_121 (
    .io_i_pj(Black_121_io_i_pj),
    .io_i_gj(Black_121_io_i_gj),
    .io_i_pk(Black_121_io_i_pk),
    .io_i_gk(Black_121_io_i_gk),
    .io_o_g(Black_121_io_o_g),
    .io_o_p(Black_121_io_o_p)
  );

  wire  PG_122_io_i_a;
  wire  PG_122_io_i_b;
  wire  PG_122_io_o_p;
  wire  PG_122_io_o_g;
  PG PG_122 (
    .io_i_a(PG_122_io_i_a),
    .io_i_b(PG_122_io_i_b),
    .io_o_p(PG_122_io_o_p),
    .io_o_g(PG_122_io_o_g)
  );

  wire  Black_123_io_i_pj;
  wire  Black_123_io_i_gj;
  wire  Black_123_io_i_pk;
  wire  Black_123_io_i_gk;
  wire  Black_123_io_o_g;
  wire  Black_123_io_o_p;
  Black Black_123 (
    .io_i_pj(Black_123_io_i_pj),
    .io_i_gj(Black_123_io_i_gj),
    .io_i_pk(Black_123_io_i_pk),
    .io_i_gk(Black_123_io_i_gk),
    .io_o_g(Black_123_io_o_g),
    .io_o_p(Black_123_io_o_p)
  );

  wire  Black_125_io_i_pj;
  wire  Black_125_io_i_gj;
  wire  Black_125_io_i_pk;
  wire  Black_125_io_i_gk;
  wire  Black_125_io_o_g;
  wire  Black_125_io_o_p;
  Black Black_125 (
    .io_i_pj(Black_125_io_i_pj),
    .io_i_gj(Black_125_io_i_gj),
    .io_i_pk(Black_125_io_i_pk),
    .io_i_gk(Black_125_io_i_gk),
    .io_o_g(Black_125_io_o_g),
    .io_o_p(Black_125_io_o_p)
  );

  wire  Black_127_io_i_pj;
  wire  Black_127_io_i_gj;
  wire  Black_127_io_i_pk;
  wire  Black_127_io_i_gk;
  wire  Black_127_io_o_g;
  wire  Black_127_io_o_p;
  Black Black_127 (
    .io_i_pj(Black_127_io_i_pj),
    .io_i_gj(Black_127_io_i_gj),
    .io_i_pk(Black_127_io_i_pk),
    .io_i_gk(Black_127_io_i_gk),
    .io_o_g(Black_127_io_o_g),
    .io_o_p(Black_127_io_o_p)
  );

  wire  Black_133_io_i_pj;
  wire  Black_133_io_i_gj;
  wire  Black_133_io_i_pk;
  wire  Black_133_io_i_gk;
  wire  Black_133_io_o_g;
  wire  Black_133_io_o_p;
  Black Black_133 (
    .io_i_pj(Black_133_io_i_pj),
    .io_i_gj(Black_133_io_i_gj),
    .io_i_pk(Black_133_io_i_pk),
    .io_i_gk(Black_133_io_i_gk),
    .io_o_g(Black_133_io_o_g),
    .io_o_p(Black_133_io_o_p)
  );

  wire  Black_135_io_i_pj;
  wire  Black_135_io_i_gj;
  wire  Black_135_io_i_pk;
  wire  Black_135_io_i_gk;
  wire  Black_135_io_o_g;
  wire  Black_135_io_o_p;
  Black Black_135 (
    .io_i_pj(Black_135_io_i_pj),
    .io_i_gj(Black_135_io_i_gj),
    .io_i_pk(Black_135_io_i_pk),
    .io_i_gk(Black_135_io_i_gk),
    .io_o_g(Black_135_io_o_g),
    .io_o_p(Black_135_io_o_p)
  );

  wire  Black_145_io_i_pj;
  wire  Black_145_io_i_gj;
  wire  Black_145_io_i_pk;
  wire  Black_145_io_i_gk;
  wire  Black_145_io_o_g;
  wire  Black_145_io_o_p;
  Black Black_145 (
    .io_i_pj(Black_145_io_i_pj),
    .io_i_gj(Black_145_io_i_gj),
    .io_i_pk(Black_145_io_i_pk),
    .io_i_gk(Black_145_io_i_gk),
    .io_o_g(Black_145_io_o_g),
    .io_o_p(Black_145_io_o_p)
  );

  wire  Black_149_io_i_pj;
  wire  Black_149_io_i_gj;
  wire  Black_149_io_i_pk;
  wire  Black_149_io_i_gk;
  wire  Black_149_io_o_g;
  wire  Black_149_io_o_p;
  Black Black_149 (
    .io_i_pj(Black_149_io_i_pj),
    .io_i_gj(Black_149_io_i_gj),
    .io_i_pk(Black_149_io_i_pk),
    .io_i_gk(Black_149_io_i_gk),
    .io_o_g(Black_149_io_o_g),
    .io_o_p(Black_149_io_o_p)
  );

  wire  PG_150_io_i_a;
  wire  PG_150_io_i_b;
  wire  PG_150_io_o_p;
  wire  PG_150_io_o_g;
  PG PG_150 (
    .io_i_a(PG_150_io_i_a),
    .io_i_b(PG_150_io_i_b),
    .io_o_p(PG_150_io_o_p),
    .io_o_g(PG_150_io_o_g)
  );

  wire  Black_152_io_i_pj;
  wire  Black_152_io_i_gj;
  wire  Black_152_io_i_pk;
  wire  Black_152_io_i_gk;
  wire  Black_152_io_o_g;
  wire  Black_152_io_o_p;
  Black Black_152 (
    .io_i_pj(Black_152_io_i_pj),
    .io_i_gj(Black_152_io_i_gj),
    .io_i_pk(Black_152_io_i_pk),
    .io_i_gk(Black_152_io_i_gk),
    .io_o_g(Black_152_io_o_g),
    .io_o_p(Black_152_io_o_p)
  );

  wire  Black_153_io_i_pj;
  wire  Black_153_io_i_gj;
  wire  Black_153_io_i_pk;
  wire  Black_153_io_i_gk;
  wire  Black_153_io_o_g;
  wire  Black_153_io_o_p;
  Black Black_153 (
    .io_i_pj(Black_153_io_i_pj),
    .io_i_gj(Black_153_io_i_gj),
    .io_i_pk(Black_153_io_i_pk),
    .io_i_gk(Black_153_io_i_gk),
    .io_o_g(Black_153_io_o_g),
    .io_o_p(Black_153_io_o_p)
  );

  wire  Black_160_io_i_pj;
  wire  Black_160_io_i_gj;
  wire  Black_160_io_i_pk;
  wire  Black_160_io_i_gk;
  wire  Black_160_io_o_g;
  wire  Black_160_io_o_p;
  Black Black_160 (
    .io_i_pj(Black_160_io_i_pj),
    .io_i_gj(Black_160_io_i_gj),
    .io_i_pk(Black_160_io_i_pk),
    .io_i_gk(Black_160_io_i_gk),
    .io_o_g(Black_160_io_o_g),
    .io_o_p(Black_160_io_o_p)
  );

  wire  Black_162_io_i_pj;
  wire  Black_162_io_i_gj;
  wire  Black_162_io_i_pk;
  wire  Black_162_io_i_gk;
  wire  Black_162_io_o_g;
  wire  Black_162_io_o_p;
  Black Black_162 (
    .io_i_pj(Black_162_io_i_pj),
    .io_i_gj(Black_162_io_i_gj),
    .io_i_pk(Black_162_io_i_pk),
    .io_i_gk(Black_162_io_i_gk),
    .io_o_g(Black_162_io_o_g),
    .io_o_p(Black_162_io_o_p)
  );

  wire  Black_176_io_i_pj;
  wire  Black_176_io_i_gj;
  wire  Black_176_io_i_pk;
  wire  Black_176_io_i_gk;
  wire  Black_176_io_o_g;
  wire  Black_176_io_o_p;
  Black Black_176 (
    .io_i_pj(Black_176_io_i_pj),
    .io_i_gj(Black_176_io_i_gj),
    .io_i_pk(Black_176_io_i_pk),
    .io_i_gk(Black_176_io_i_gk),
    .io_o_g(Black_176_io_o_g),
    .io_o_p(Black_176_io_o_p)
  );

  wire  PG_177_io_i_a;
  wire  PG_177_io_i_b;
  wire  PG_177_io_o_p;
  wire  PG_177_io_o_g;
  PG PG_177 (
    .io_i_a(PG_177_io_i_a),
    .io_i_b(PG_177_io_i_b),
    .io_o_p(PG_177_io_o_p),
    .io_o_g(PG_177_io_o_g)
  );

  wire  Black_178_io_i_pj;
  wire  Black_178_io_i_gj;
  wire  Black_178_io_i_pk;
  wire  Black_178_io_i_gk;
  wire  Black_178_io_o_g;
  wire  Black_178_io_o_p;
  Black Black_178 (
    .io_i_pj(Black_178_io_i_pj),
    .io_i_gj(Black_178_io_i_gj),
    .io_i_pk(Black_178_io_i_pk),
    .io_i_gk(Black_178_io_i_gk),
    .io_o_g(Black_178_io_o_g),
    .io_o_p(Black_178_io_o_p)
  );

  wire  Black_180_io_i_pj;
  wire  Black_180_io_i_gj;
  wire  Black_180_io_i_pk;
  wire  Black_180_io_i_gk;
  wire  Black_180_io_o_g;
  wire  Black_180_io_o_p;
  Black Black_180 (
    .io_i_pj(Black_180_io_i_pj),
    .io_i_gj(Black_180_io_i_gj),
    .io_i_pk(Black_180_io_i_pk),
    .io_i_gk(Black_180_io_i_gk),
    .io_o_g(Black_180_io_o_g),
    .io_o_p(Black_180_io_o_p)
  );

  wire  Black_202_io_i_pj;
  wire  Black_202_io_i_gj;
  wire  Black_202_io_i_pk;
  wire  Black_202_io_i_gk;
  wire  Black_202_io_o_g;
  wire  Black_202_io_o_p;
  Black Black_202 (
    .io_i_pj(Black_202_io_i_pj),
    .io_i_gj(Black_202_io_i_gj),
    .io_i_pk(Black_202_io_i_pk),
    .io_i_gk(Black_202_io_i_gk),
    .io_o_g(Black_202_io_o_g),
    .io_o_p(Black_202_io_o_p)
  );

  wire  PG_203_io_i_a;
  wire  PG_203_io_i_b;
  wire  PG_203_io_o_p;
  wire  PG_203_io_o_g;
  PG PG_203 (
    .io_i_a(PG_203_io_i_a),
    .io_i_b(PG_203_io_i_b),
    .io_o_p(PG_203_io_o_p),
    .io_o_g(PG_203_io_o_g)
  );

  wire  Black_211_io_i_pj;
  wire  Black_211_io_i_gj;
  wire  Black_211_io_i_pk;
  wire  Black_211_io_i_gk;
  wire  Black_211_io_o_g;
  wire  Black_211_io_o_p;
  Black Black_211 (
    .io_i_pj(Black_211_io_i_pj),
    .io_i_gj(Black_211_io_i_gj),
    .io_i_pk(Black_211_io_i_pk),
    .io_i_gk(Black_211_io_i_gk),
    .io_o_g(Black_211_io_o_g),
    .io_o_p(Black_211_io_o_p)
  );

  wire  Black_227_io_i_pj;
  wire  Black_227_io_i_gj;
  wire  Black_227_io_i_pk;
  wire  Black_227_io_i_gk;
  wire  Black_227_io_o_g;
  wire  Black_227_io_o_p;
  Black Black_227 (
    .io_i_pj(Black_227_io_i_pj),
    .io_i_gj(Black_227_io_i_gj),
    .io_i_pk(Black_227_io_i_pk),
    .io_i_gk(Black_227_io_i_gk),
    .io_o_g(Black_227_io_o_g),
    .io_o_p(Black_227_io_o_p)
  );

  wire  PG_228_io_i_a;
  wire  PG_228_io_i_b;
  wire  PG_228_io_o_p;
  wire  PG_228_io_o_g;
  PG PG_228 (
    .io_i_a(PG_228_io_i_a),
    .io_i_b(PG_228_io_i_b),
    .io_o_p(PG_228_io_o_p),
    .io_o_g(PG_228_io_o_g)
  );

  wire  Black_229_io_i_pj;
  wire  Black_229_io_i_gj;
  wire  Black_229_io_i_pk;
  wire  Black_229_io_i_gk;
  wire  Black_229_io_o_g;
  wire  Black_229_io_o_p;
  Black Black_229 (
    .io_i_pj(Black_229_io_i_pj),
    .io_i_gj(Black_229_io_i_gj),
    .io_i_pk(Black_229_io_i_pk),
    .io_i_gk(Black_229_io_i_gk),
    .io_o_g(Black_229_io_o_g),
    .io_o_p(Black_229_io_o_p)
  );

  wire  Black_231_io_i_pj;
  wire  Black_231_io_i_gj;
  wire  Black_231_io_i_pk;
  wire  Black_231_io_i_gk;
  wire  Black_231_io_o_g;
  wire  Black_231_io_o_p;
  Black Black_231 (
    .io_i_pj(Black_231_io_i_pj),
    .io_i_gj(Black_231_io_i_gj),
    .io_i_pk(Black_231_io_i_pk),
    .io_i_gk(Black_231_io_i_gk),
    .io_o_g(Black_231_io_o_g),
    .io_o_p(Black_231_io_o_p)
  );

  wire  Black_235_io_i_pj;
  wire  Black_235_io_i_gj;
  wire  Black_235_io_i_pk;
  wire  Black_235_io_i_gk;
  wire  Black_235_io_o_g;
  wire  Black_235_io_o_p;
  Black Black_235 (
    .io_i_pj(Black_235_io_i_pj),
    .io_i_gj(Black_235_io_i_gj),
    .io_i_pk(Black_235_io_i_pk),
    .io_i_gk(Black_235_io_i_gk),
    .io_o_g(Black_235_io_o_g),
    .io_o_p(Black_235_io_o_p)
  );

  wire  Black_238_io_i_pj;
  wire  Black_238_io_i_gj;
  wire  Black_238_io_i_pk;
  wire  Black_238_io_i_gk;
  wire  Black_238_io_o_g;
  wire  Black_238_io_o_p;
  Black Black_238 (
    .io_i_pj(Black_238_io_i_pj),
    .io_i_gj(Black_238_io_i_gj),
    .io_i_pk(Black_238_io_i_pk),
    .io_i_gk(Black_238_io_i_gk),
    .io_o_g(Black_238_io_o_g),
    .io_o_p(Black_238_io_o_p)
  );

  wire  Black_240_io_i_pj;
  wire  Black_240_io_i_gj;
  wire  Black_240_io_i_pk;
  wire  Black_240_io_i_gk;
  wire  Black_240_io_o_g;
  wire  Black_240_io_o_p;
  Black Black_240 (
    .io_i_pj(Black_240_io_i_pj),
    .io_i_gj(Black_240_io_i_gj),
    .io_i_pk(Black_240_io_i_pk),
    .io_i_gk(Black_240_io_i_gk),
    .io_o_g(Black_240_io_o_g),
    .io_o_p(Black_240_io_o_p)
  );

  wire  Black_242_io_i_pj;
  wire  Black_242_io_i_gj;
  wire  Black_242_io_i_pk;
  wire  Black_242_io_i_gk;
  wire  Black_242_io_o_g;
  wire  Black_242_io_o_p;
  Black Black_242 (
    .io_i_pj(Black_242_io_i_pj),
    .io_i_gj(Black_242_io_i_gj),
    .io_i_pk(Black_242_io_i_pk),
    .io_i_gk(Black_242_io_i_gk),
    .io_o_g(Black_242_io_o_g),
    .io_o_p(Black_242_io_o_p)
  );

  wire  Black_246_io_i_pj;
  wire  Black_246_io_i_gj;
  wire  Black_246_io_i_pk;
  wire  Black_246_io_i_gk;
  wire  Black_246_io_o_g;
  wire  Black_246_io_o_p;
  Black Black_246 (
    .io_i_pj(Black_246_io_i_pj),
    .io_i_gj(Black_246_io_i_gj),
    .io_i_pk(Black_246_io_i_pk),
    .io_i_gk(Black_246_io_i_gk),
    .io_o_g(Black_246_io_o_g),
    .io_o_p(Black_246_io_o_p)
  );

  wire  Black_248_io_i_pj;
  wire  Black_248_io_i_gj;
  wire  Black_248_io_i_pk;
  wire  Black_248_io_i_gk;
  wire  Black_248_io_o_g;
  wire  Black_248_io_o_p;
  Black Black_248 (
    .io_i_pj(Black_248_io_i_pj),
    .io_i_gj(Black_248_io_i_gj),
    .io_i_pk(Black_248_io_i_pk),
    .io_i_gk(Black_248_io_i_gk),
    .io_o_g(Black_248_io_o_g),
    .io_o_p(Black_248_io_o_p)
  );

  wire  Black_251_io_i_pj;
  wire  Black_251_io_i_gj;
  wire  Black_251_io_i_pk;
  wire  Black_251_io_i_gk;
  wire  Black_251_io_o_g;
  wire  Black_251_io_o_p;
  Black Black_251 (
    .io_i_pj(Black_251_io_i_pj),
    .io_i_gj(Black_251_io_i_gj),
    .io_i_pk(Black_251_io_i_pk),
    .io_i_gk(Black_251_io_i_gk),
    .io_o_g(Black_251_io_o_g),
    .io_o_p(Black_251_io_o_p)
  );

  wire  PG_252_io_i_a;
  wire  PG_252_io_i_b;
  wire  PG_252_io_o_p;
  wire  PG_252_io_o_g;
  PG PG_252 (
    .io_i_a(PG_252_io_i_a),
    .io_i_b(PG_252_io_i_b),
    .io_o_p(PG_252_io_o_p),
    .io_o_g(PG_252_io_o_g)
  );

  wire  Black_253_io_i_pj;
  wire  Black_253_io_i_gj;
  wire  Black_253_io_i_pk;
  wire  Black_253_io_i_gk;
  wire  Black_253_io_o_g;
  wire  Black_253_io_o_p;
  Black Black_253 (
    .io_i_pj(Black_253_io_i_pj),
    .io_i_gj(Black_253_io_i_gj),
    .io_i_pk(Black_253_io_i_pk),
    .io_i_gk(Black_253_io_i_gk),
    .io_o_g(Black_253_io_o_g),
    .io_o_p(Black_253_io_o_p)
  );

  wire  Black_254_io_i_pj;
  wire  Black_254_io_i_gj;
  wire  Black_254_io_i_pk;
  wire  Black_254_io_i_gk;
  wire  Black_254_io_o_g;
  wire  Black_254_io_o_p;
  Black Black_254 (
    .io_i_pj(Black_254_io_i_pj),
    .io_i_gj(Black_254_io_i_gj),
    .io_i_pk(Black_254_io_i_pk),
    .io_i_gk(Black_254_io_i_gk),
    .io_o_g(Black_254_io_o_g),
    .io_o_p(Black_254_io_o_p)
  );

  wire  Black_257_io_i_pj;
  wire  Black_257_io_i_gj;
  wire  Black_257_io_i_pk;
  wire  Black_257_io_i_gk;
  wire  Black_257_io_o_g;
  wire  Black_257_io_o_p;
  Black Black_257 (
    .io_i_pj(Black_257_io_i_pj),
    .io_i_gj(Black_257_io_i_gj),
    .io_i_pk(Black_257_io_i_pk),
    .io_i_gk(Black_257_io_i_gk),
    .io_o_g(Black_257_io_o_g),
    .io_o_p(Black_257_io_o_p)
  );

  wire  Black_258_io_i_pj;
  wire  Black_258_io_i_gj;
  wire  Black_258_io_i_pk;
  wire  Black_258_io_i_gk;
  wire  Black_258_io_o_g;
  wire  Black_258_io_o_p;
  Black Black_258 (
    .io_i_pj(Black_258_io_i_pj),
    .io_i_gj(Black_258_io_i_gj),
    .io_i_pk(Black_258_io_i_pk),
    .io_i_gk(Black_258_io_i_gk),
    .io_o_g(Black_258_io_o_g),
    .io_o_p(Black_258_io_o_p)
  );

  wire  Black_263_io_i_pj;
  wire  Black_263_io_i_gj;
  wire  Black_263_io_i_pk;
  wire  Black_263_io_i_gk;
  wire  Black_263_io_o_g;
  wire  Black_263_io_o_p;
  Black Black_263 (
    .io_i_pj(Black_263_io_i_pj),
    .io_i_gj(Black_263_io_i_gj),
    .io_i_pk(Black_263_io_i_pk),
    .io_i_gk(Black_263_io_i_gk),
    .io_o_g(Black_263_io_o_g),
    .io_o_p(Black_263_io_o_p)
  );

  wire  Black_274_io_i_pj;
  wire  Black_274_io_i_gj;
  wire  Black_274_io_i_pk;
  wire  Black_274_io_i_gk;
  wire  Black_274_io_o_g;
  wire  Black_274_io_o_p;
  Black Black_274 (
    .io_i_pj(Black_274_io_i_pj),
    .io_i_gj(Black_274_io_i_gj),
    .io_i_pk(Black_274_io_i_pk),
    .io_i_gk(Black_274_io_i_gk),
    .io_o_g(Black_274_io_o_g),
    .io_o_p(Black_274_io_o_p)
  );

  wire  PG_275_io_i_a;
  wire  PG_275_io_i_b;
  wire  PG_275_io_o_p;
  wire  PG_275_io_o_g;
  PG PG_275 (
    .io_i_a(PG_275_io_i_a),
    .io_i_b(PG_275_io_i_b),
    .io_o_p(PG_275_io_o_p),
    .io_o_g(PG_275_io_o_g)
  );

  wire  Black_276_io_i_pj;
  wire  Black_276_io_i_gj;
  wire  Black_276_io_i_pk;
  wire  Black_276_io_i_gk;
  wire  Black_276_io_o_g;
  wire  Black_276_io_o_p;
  Black Black_276 (
    .io_i_pj(Black_276_io_i_pj),
    .io_i_gj(Black_276_io_i_gj),
    .io_i_pk(Black_276_io_i_pk),
    .io_i_gk(Black_276_io_i_gk),
    .io_o_g(Black_276_io_o_g),
    .io_o_p(Black_276_io_o_p)
  );

  wire  Black_280_io_i_pj;
  wire  Black_280_io_i_gj;
  wire  Black_280_io_i_pk;
  wire  Black_280_io_i_gk;
  wire  Black_280_io_o_g;
  wire  Black_280_io_o_p;
  Black Black_280 (
    .io_i_pj(Black_280_io_i_pj),
    .io_i_gj(Black_280_io_i_gj),
    .io_i_pk(Black_280_io_i_pk),
    .io_i_gk(Black_280_io_i_gk),
    .io_o_g(Black_280_io_o_g),
    .io_o_p(Black_280_io_o_p)
  );

  wire  Black_289_io_i_pj;
  wire  Black_289_io_i_gj;
  wire  Black_289_io_i_pk;
  wire  Black_289_io_i_gk;
  wire  Black_289_io_o_g;
  wire  Black_289_io_o_p;
  Black Black_289 (
    .io_i_pj(Black_289_io_i_pj),
    .io_i_gj(Black_289_io_i_gj),
    .io_i_pk(Black_289_io_i_pk),
    .io_i_gk(Black_289_io_i_gk),
    .io_o_g(Black_289_io_o_g),
    .io_o_p(Black_289_io_o_p)
  );

  wire  Black_296_io_i_pj;
  wire  Black_296_io_i_gj;
  wire  Black_296_io_i_pk;
  wire  Black_296_io_i_gk;
  wire  Black_296_io_o_g;
  wire  Black_296_io_o_p;
  Black Black_296 (
    .io_i_pj(Black_296_io_i_pj),
    .io_i_gj(Black_296_io_i_gj),
    .io_i_pk(Black_296_io_i_pk),
    .io_i_gk(Black_296_io_i_gk),
    .io_o_g(Black_296_io_o_g),
    .io_o_p(Black_296_io_o_p)
  );

  wire  PG_297_io_i_a;
  wire  PG_297_io_i_b;
  wire  PG_297_io_o_p;
  wire  PG_297_io_o_g;
  PG PG_297 (
    .io_i_a(PG_297_io_i_a),
    .io_i_b(PG_297_io_i_b),
    .io_o_p(PG_297_io_o_p),
    .io_o_g(PG_297_io_o_g)
  );

  wire  Black_298_io_i_pj;
  wire  Black_298_io_i_gj;
  wire  Black_298_io_i_pk;
  wire  Black_298_io_i_gk;
  wire  Black_298_io_o_g;
  wire  Black_298_io_o_p;
  Black Black_298 (
    .io_i_pj(Black_298_io_i_pj),
    .io_i_gj(Black_298_io_i_gj),
    .io_i_pk(Black_298_io_i_pk),
    .io_i_gk(Black_298_io_i_gk),
    .io_o_g(Black_298_io_o_g),
    .io_o_p(Black_298_io_o_p)
  );

  wire  Black_317_io_i_pj;
  wire  Black_317_io_i_gj;
  wire  Black_317_io_i_pk;
  wire  Black_317_io_i_gk;
  wire  Black_317_io_o_g;
  wire  Black_317_io_o_p;
  Black Black_317 (
    .io_i_pj(Black_317_io_i_pj),
    .io_i_gj(Black_317_io_i_gj),
    .io_i_pk(Black_317_io_i_pk),
    .io_i_gk(Black_317_io_i_gk),
    .io_o_g(Black_317_io_o_g),
    .io_o_p(Black_317_io_o_p)
  );

  wire  PG_318_io_i_a;
  wire  PG_318_io_i_b;
  wire  PG_318_io_o_p;
  wire  PG_318_io_o_g;
  PG PG_318 (
    .io_i_a(PG_318_io_i_a),
    .io_i_b(PG_318_io_i_b),
    .io_o_p(PG_318_io_o_p),
    .io_o_g(PG_318_io_o_g)
  );

  wire  Black_319_io_i_pj;
  wire  Black_319_io_i_gj;
  wire  Black_319_io_i_pk;
  wire  Black_319_io_i_gk;
  wire  Black_319_io_o_g;
  wire  Black_319_io_o_p;
  Black Black_319 (
    .io_i_pj(Black_319_io_i_pj),
    .io_i_gj(Black_319_io_i_gj),
    .io_i_pk(Black_319_io_i_pk),
    .io_i_gk(Black_319_io_i_gk),
    .io_o_g(Black_319_io_o_g),
    .io_o_p(Black_319_io_o_p)
  );

  wire  Black_320_io_i_pj;
  wire  Black_320_io_i_gj;
  wire  Black_320_io_i_pk;
  wire  Black_320_io_i_gk;
  wire  Black_320_io_o_g;
  wire  Black_320_io_o_p;
  Black Black_320 (
    .io_i_pj(Black_320_io_i_pj),
    .io_i_gj(Black_320_io_i_gj),
    .io_i_pk(Black_320_io_i_pk),
    .io_i_gk(Black_320_io_i_gk),
    .io_o_g(Black_320_io_o_g),
    .io_o_p(Black_320_io_o_p)
  );

  wire  Black_321_io_i_pj;
  wire  Black_321_io_i_gj;
  wire  Black_321_io_i_pk;
  wire  Black_321_io_i_gk;
  wire  Black_321_io_o_g;
  wire  Black_321_io_o_p;
  Black Black_321 (
    .io_i_pj(Black_321_io_i_pj),
    .io_i_gj(Black_321_io_i_gj),
    .io_i_pk(Black_321_io_i_pk),
    .io_i_gk(Black_321_io_i_gk),
    .io_o_g(Black_321_io_o_g),
    .io_o_p(Black_321_io_o_p)
  );

  wire  Black_337_io_i_pj;
  wire  Black_337_io_i_gj;
  wire  Black_337_io_i_pk;
  wire  Black_337_io_i_gk;
  wire  Black_337_io_o_g;
  wire  Black_337_io_o_p;
  Black Black_337 (
    .io_i_pj(Black_337_io_i_pj),
    .io_i_gj(Black_337_io_i_gj),
    .io_i_pk(Black_337_io_i_pk),
    .io_i_gk(Black_337_io_i_gk),
    .io_o_g(Black_337_io_o_g),
    .io_o_p(Black_337_io_o_p)
  );

  wire  PG_338_io_i_a;
  wire  PG_338_io_i_b;
  wire  PG_338_io_o_p;
  wire  PG_338_io_o_g;
  PG PG_338 (
    .io_i_a(PG_338_io_i_a),
    .io_i_b(PG_338_io_i_b),
    .io_o_p(PG_338_io_o_p),
    .io_o_g(PG_338_io_o_g)
  );

  wire  Black_340_io_i_pj;
  wire  Black_340_io_i_gj;
  wire  Black_340_io_i_pk;
  wire  Black_340_io_i_gk;
  wire  Black_340_io_o_g;
  wire  Black_340_io_o_p;
  Black Black_340 (
    .io_i_pj(Black_340_io_i_pj),
    .io_i_gj(Black_340_io_i_gj),
    .io_i_pk(Black_340_io_i_pk),
    .io_i_gk(Black_340_io_i_gk),
    .io_o_g(Black_340_io_o_g),
    .io_o_p(Black_340_io_o_p)
  );

  wire  Black_352_io_i_pj;
  wire  Black_352_io_i_gj;
  wire  Black_352_io_i_pk;
  wire  Black_352_io_i_gk;
  wire  Black_352_io_o_g;
  wire  Black_352_io_o_p;
  Black Black_352 (
    .io_i_pj(Black_352_io_i_pj),
    .io_i_gj(Black_352_io_i_gj),
    .io_i_pk(Black_352_io_i_pk),
    .io_i_gk(Black_352_io_i_gk),
    .io_o_g(Black_352_io_o_g),
    .io_o_p(Black_352_io_o_p)
  );

  wire  Black_356_io_i_pj;
  wire  Black_356_io_i_gj;
  wire  Black_356_io_i_pk;
  wire  Black_356_io_i_gk;
  wire  Black_356_io_o_g;
  wire  Black_356_io_o_p;
  Black Black_356 (
    .io_i_pj(Black_356_io_i_pj),
    .io_i_gj(Black_356_io_i_gj),
    .io_i_pk(Black_356_io_i_pk),
    .io_i_gk(Black_356_io_i_gk),
    .io_o_g(Black_356_io_o_g),
    .io_o_p(Black_356_io_o_p)
  );

  wire  PG_357_io_i_a;
  wire  PG_357_io_i_b;
  wire  PG_357_io_o_p;
  wire  PG_357_io_o_g;
  PG PG_357 (
    .io_i_a(PG_357_io_i_a),
    .io_i_b(PG_357_io_i_b),
    .io_o_p(PG_357_io_o_p),
    .io_o_g(PG_357_io_o_g)
  );

  wire  Black_358_io_i_pj;
  wire  Black_358_io_i_gj;
  wire  Black_358_io_i_pk;
  wire  Black_358_io_i_gk;
  wire  Black_358_io_o_g;
  wire  Black_358_io_o_p;
  Black Black_358 (
    .io_i_pj(Black_358_io_i_pj),
    .io_i_gj(Black_358_io_i_gj),
    .io_i_pk(Black_358_io_i_pk),
    .io_i_gk(Black_358_io_i_gk),
    .io_o_g(Black_358_io_o_g),
    .io_o_p(Black_358_io_o_p)
  );

  wire  Black_363_io_i_pj;
  wire  Black_363_io_i_gj;
  wire  Black_363_io_i_pk;
  wire  Black_363_io_i_gk;
  wire  Black_363_io_o_g;
  wire  Black_363_io_o_p;
  Black Black_363 (
    .io_i_pj(Black_363_io_i_pj),
    .io_i_gj(Black_363_io_i_gj),
    .io_i_pk(Black_363_io_i_pk),
    .io_i_gk(Black_363_io_i_gk),
    .io_o_g(Black_363_io_o_g),
    .io_o_p(Black_363_io_o_p)
  );

  wire  Black_374_io_i_pj;
  wire  Black_374_io_i_gj;
  wire  Black_374_io_i_pk;
  wire  Black_374_io_i_gk;
  wire  Black_374_io_o_g;
  wire  Black_374_io_o_p;
  Black Black_374 (
    .io_i_pj(Black_374_io_i_pj),
    .io_i_gj(Black_374_io_i_gj),
    .io_i_pk(Black_374_io_i_pk),
    .io_i_gk(Black_374_io_i_gk),
    .io_o_g(Black_374_io_o_g),
    .io_o_p(Black_374_io_o_p)
  );

  wire  PG_375_io_i_a;
  wire  PG_375_io_i_b;
  wire  PG_375_io_o_p;
  wire  PG_375_io_o_g;
  PG PG_375 (
    .io_i_a(PG_375_io_i_a),
    .io_i_b(PG_375_io_i_b),
    .io_o_p(PG_375_io_o_p),
    .io_o_g(PG_375_io_o_g)
  );

  wire  Black_391_io_i_pj;
  wire  Black_391_io_i_gj;
  wire  Black_391_io_i_pk;
  wire  Black_391_io_i_gk;
  wire  Black_391_io_o_g;
  wire  Black_391_io_o_p;
  Black Black_391 (
    .io_i_pj(Black_391_io_i_pj),
    .io_i_gj(Black_391_io_i_gj),
    .io_i_pk(Black_391_io_i_pk),
    .io_i_gk(Black_391_io_i_gk),
    .io_o_g(Black_391_io_o_g),
    .io_o_p(Black_391_io_o_p)
  );

  wire  PG_392_io_i_a;
  wire  PG_392_io_i_b;
  wire  PG_392_io_o_p;
  wire  PG_392_io_o_g;
  PG PG_392 (
    .io_i_a(PG_392_io_i_a),
    .io_i_b(PG_392_io_i_b),
    .io_o_p(PG_392_io_o_p),
    .io_o_g(PG_392_io_o_g)
  );

  wire  Black_393_io_i_pj;
  wire  Black_393_io_i_gj;
  wire  Black_393_io_i_pk;
  wire  Black_393_io_i_gk;
  wire  Black_393_io_o_g;
  wire  Black_393_io_o_p;
  Black Black_393 (
    .io_i_pj(Black_393_io_i_pj),
    .io_i_gj(Black_393_io_i_gj),
    .io_i_pk(Black_393_io_i_pk),
    .io_i_gk(Black_393_io_i_gk),
    .io_o_g(Black_393_io_o_g),
    .io_o_p(Black_393_io_o_p)
  );

  wire  Black_394_io_i_pj;
  wire  Black_394_io_i_gj;
  wire  Black_394_io_i_pk;
  wire  Black_394_io_i_gk;
  wire  Black_394_io_o_g;
  wire  Black_394_io_o_p;
  Black Black_394 (
    .io_i_pj(Black_394_io_i_pj),
    .io_i_gj(Black_394_io_i_gj),
    .io_i_pk(Black_394_io_i_pk),
    .io_i_gk(Black_394_io_i_gk),
    .io_o_g(Black_394_io_o_g),
    .io_o_p(Black_394_io_o_p)
  );

  wire  Black_395_io_i_pj;
  wire  Black_395_io_i_gj;
  wire  Black_395_io_i_pk;
  wire  Black_395_io_i_gk;
  wire  Black_395_io_o_g;
  wire  Black_395_io_o_p;
  Black Black_395 (
    .io_i_pj(Black_395_io_i_pj),
    .io_i_gj(Black_395_io_i_gj),
    .io_i_pk(Black_395_io_i_pk),
    .io_i_gk(Black_395_io_i_gk),
    .io_o_g(Black_395_io_o_g),
    .io_o_p(Black_395_io_o_p)
  );

  wire  Black_396_io_i_pj;
  wire  Black_396_io_i_gj;
  wire  Black_396_io_i_pk;
  wire  Black_396_io_i_gk;
  wire  Black_396_io_o_g;
  wire  Black_396_io_o_p;
  Black Black_396 (
    .io_i_pj(Black_396_io_i_pj),
    .io_i_gj(Black_396_io_i_gj),
    .io_i_pk(Black_396_io_i_pk),
    .io_i_gk(Black_396_io_i_gk),
    .io_o_g(Black_396_io_o_g),
    .io_o_p(Black_396_io_o_p)
  );

  wire  Black_398_io_i_pj;
  wire  Black_398_io_i_gj;
  wire  Black_398_io_i_pk;
  wire  Black_398_io_i_gk;
  wire  Black_398_io_o_g;
  wire  Black_398_io_o_p;
  Black Black_398 (
    .io_i_pj(Black_398_io_i_pj),
    .io_i_gj(Black_398_io_i_gj),
    .io_i_pk(Black_398_io_i_pk),
    .io_i_gk(Black_398_io_i_gk),
    .io_o_g(Black_398_io_o_g),
    .io_o_p(Black_398_io_o_p)
  );

  wire  Black_399_io_i_pj;
  wire  Black_399_io_i_gj;
  wire  Black_399_io_i_pk;
  wire  Black_399_io_i_gk;
  wire  Black_399_io_o_g;
  wire  Black_399_io_o_p;
  Black Black_399 (
    .io_i_pj(Black_399_io_i_pj),
    .io_i_gj(Black_399_io_i_gj),
    .io_i_pk(Black_399_io_i_pk),
    .io_i_gk(Black_399_io_i_gk),
    .io_o_g(Black_399_io_o_g),
    .io_o_p(Black_399_io_o_p)
  );

  wire  Black_400_io_i_pj;
  wire  Black_400_io_i_gj;
  wire  Black_400_io_i_pk;
  wire  Black_400_io_i_gk;
  wire  Black_400_io_o_g;
  wire  Black_400_io_o_p;
  Black Black_400 (
    .io_i_pj(Black_400_io_i_pj),
    .io_i_gj(Black_400_io_i_gj),
    .io_i_pk(Black_400_io_i_pk),
    .io_i_gk(Black_400_io_i_gk),
    .io_o_g(Black_400_io_o_g),
    .io_o_p(Black_400_io_o_p)
  );

  wire  Black_403_io_i_pj;
  wire  Black_403_io_i_gj;
  wire  Black_403_io_i_pk;
  wire  Black_403_io_i_gk;
  wire  Black_403_io_o_g;
  wire  Black_403_io_o_p;
  Black Black_403 (
    .io_i_pj(Black_403_io_i_pj),
    .io_i_gj(Black_403_io_i_gj),
    .io_i_pk(Black_403_io_i_pk),
    .io_i_gk(Black_403_io_i_gk),
    .io_o_g(Black_403_io_o_g),
    .io_o_p(Black_403_io_o_p)
  );

  wire  Black_407_io_i_pj;
  wire  Black_407_io_i_gj;
  wire  Black_407_io_i_pk;
  wire  Black_407_io_i_gk;
  wire  Black_407_io_o_g;
  wire  Black_407_io_o_p;
  Black Black_407 (
    .io_i_pj(Black_407_io_i_pj),
    .io_i_gj(Black_407_io_i_gj),
    .io_i_pk(Black_407_io_i_pk),
    .io_i_gk(Black_407_io_i_gk),
    .io_o_g(Black_407_io_o_g),
    .io_o_p(Black_407_io_o_p)
  );

  wire  PG_408_io_i_a;
  wire  PG_408_io_i_b;
  wire  PG_408_io_o_p;
  wire  PG_408_io_o_g;
  PG PG_408 (
    .io_i_a(PG_408_io_i_a),
    .io_i_b(PG_408_io_i_b),
    .io_o_p(PG_408_io_o_p),
    .io_o_g(PG_408_io_o_g)
  );

  wire  Black_414_io_i_pj;
  wire  Black_414_io_i_gj;
  wire  Black_414_io_i_pk;
  wire  Black_414_io_i_gk;
  wire  Black_414_io_o_g;
  wire  Black_414_io_o_p;
  Black Black_414 (
    .io_i_pj(Black_414_io_i_pj),
    .io_i_gj(Black_414_io_i_gj),
    .io_i_pk(Black_414_io_i_pk),
    .io_i_gk(Black_414_io_i_gk),
    .io_o_g(Black_414_io_o_g),
    .io_o_p(Black_414_io_o_p)
  );

  wire  Black_416_io_i_pj;
  wire  Black_416_io_i_gj;
  wire  Black_416_io_i_pk;
  wire  Black_416_io_i_gk;
  wire  Black_416_io_o_g;
  wire  Black_416_io_o_p;
  Black Black_416 (
    .io_i_pj(Black_416_io_i_pj),
    .io_i_gj(Black_416_io_i_gj),
    .io_i_pk(Black_416_io_i_pk),
    .io_i_gk(Black_416_io_i_gk),
    .io_o_g(Black_416_io_o_g),
    .io_o_p(Black_416_io_o_p)
  );

  wire  Black_422_io_i_pj;
  wire  Black_422_io_i_gj;
  wire  Black_422_io_i_pk;
  wire  Black_422_io_i_gk;
  wire  Black_422_io_o_g;
  wire  Black_422_io_o_p;
  Black Black_422 (
    .io_i_pj(Black_422_io_i_pj),
    .io_i_gj(Black_422_io_i_gj),
    .io_i_pk(Black_422_io_i_pk),
    .io_i_gk(Black_422_io_i_gk),
    .io_o_g(Black_422_io_o_g),
    .io_o_p(Black_422_io_o_p)
  );

  wire  PG_423_io_i_a;
  wire  PG_423_io_i_b;
  wire  PG_423_io_o_p;
  wire  PG_423_io_o_g;
  PG PG_423 (
    .io_i_a(PG_423_io_i_a),
    .io_i_b(PG_423_io_i_b),
    .io_o_p(PG_423_io_o_p),
    .io_o_g(PG_423_io_o_g)
  );

  wire  Black_428_io_i_pj;
  wire  Black_428_io_i_gj;
  wire  Black_428_io_i_pk;
  wire  Black_428_io_i_gk;
  wire  Black_428_io_o_g;
  wire  Black_428_io_o_p;
  Black Black_428 (
    .io_i_pj(Black_428_io_i_pj),
    .io_i_gj(Black_428_io_i_gj),
    .io_i_pk(Black_428_io_i_pk),
    .io_i_gk(Black_428_io_i_gk),
    .io_o_g(Black_428_io_o_g),
    .io_o_p(Black_428_io_o_p)
  );

  wire  Black_432_io_i_pj;
  wire  Black_432_io_i_gj;
  wire  Black_432_io_i_pk;
  wire  Black_432_io_i_gk;
  wire  Black_432_io_o_g;
  wire  Black_432_io_o_p;
  Black Black_432 (
    .io_i_pj(Black_432_io_i_pj),
    .io_i_gj(Black_432_io_i_gj),
    .io_i_pk(Black_432_io_i_pk),
    .io_i_gk(Black_432_io_i_gk),
    .io_o_g(Black_432_io_o_g),
    .io_o_p(Black_432_io_o_p)
  );

  wire  Black_436_io_i_pj;
  wire  Black_436_io_i_gj;
  wire  Black_436_io_i_pk;
  wire  Black_436_io_i_gk;
  wire  Black_436_io_o_g;
  wire  Black_436_io_o_p;
  Black Black_436 (
    .io_i_pj(Black_436_io_i_pj),
    .io_i_gj(Black_436_io_i_gj),
    .io_i_pk(Black_436_io_i_pk),
    .io_i_gk(Black_436_io_i_gk),
    .io_o_g(Black_436_io_o_g),
    .io_o_p(Black_436_io_o_p)
  );

  wire  PG_437_io_i_a;
  wire  PG_437_io_i_b;
  wire  PG_437_io_o_p;
  wire  PG_437_io_o_g;
  PG PG_437 (
    .io_i_a(PG_437_io_i_a),
    .io_i_b(PG_437_io_i_b),
    .io_o_p(PG_437_io_o_p),
    .io_o_g(PG_437_io_o_g)
  );

  wire  Black_438_io_i_pj;
  wire  Black_438_io_i_gj;
  wire  Black_438_io_i_pk;
  wire  Black_438_io_i_gk;
  wire  Black_438_io_o_g;
  wire  Black_438_io_o_p;
  Black Black_438 (
    .io_i_pj(Black_438_io_i_pj),
    .io_i_gj(Black_438_io_i_gj),
    .io_i_pk(Black_438_io_i_pk),
    .io_i_gk(Black_438_io_i_gk),
    .io_o_g(Black_438_io_o_g),
    .io_o_p(Black_438_io_o_p)
  );

  wire  Black_441_io_i_pj;
  wire  Black_441_io_i_gj;
  wire  Black_441_io_i_pk;
  wire  Black_441_io_i_gk;
  wire  Black_441_io_o_g;
  wire  Black_441_io_o_p;
  Black Black_441 (
    .io_i_pj(Black_441_io_i_pj),
    .io_i_gj(Black_441_io_i_gj),
    .io_i_pk(Black_441_io_i_pk),
    .io_i_gk(Black_441_io_i_gk),
    .io_o_g(Black_441_io_o_g),
    .io_o_p(Black_441_io_o_p)
  );

  wire  Black_448_io_i_pj;
  wire  Black_448_io_i_gj;
  wire  Black_448_io_i_pk;
  wire  Black_448_io_i_gk;
  wire  Black_448_io_o_g;
  wire  Black_448_io_o_p;
  Black Black_448 (
    .io_i_pj(Black_448_io_i_pj),
    .io_i_gj(Black_448_io_i_gj),
    .io_i_pk(Black_448_io_i_pk),
    .io_i_gk(Black_448_io_i_gk),
    .io_o_g(Black_448_io_o_g),
    .io_o_p(Black_448_io_o_p)
  );

  wire  Black_449_io_i_pj;
  wire  Black_449_io_i_gj;
  wire  Black_449_io_i_pk;
  wire  Black_449_io_i_gk;
  wire  Black_449_io_o_g;
  wire  Black_449_io_o_p;
  Black Black_449 (
    .io_i_pj(Black_449_io_i_pj),
    .io_i_gj(Black_449_io_i_gj),
    .io_i_pk(Black_449_io_i_pk),
    .io_i_gk(Black_449_io_i_gk),
    .io_o_g(Black_449_io_o_g),
    .io_o_p(Black_449_io_o_p)
  );

  wire  PG_450_io_i_a;
  wire  PG_450_io_i_b;
  wire  PG_450_io_o_p;
  wire  PG_450_io_o_g;
  PG PG_450 (
    .io_i_a(PG_450_io_i_a),
    .io_i_b(PG_450_io_i_b),
    .io_o_p(PG_450_io_o_p),
    .io_o_g(PG_450_io_o_g)
  );

  wire  Black_451_io_i_pj;
  wire  Black_451_io_i_gj;
  wire  Black_451_io_i_pk;
  wire  Black_451_io_i_gk;
  wire  Black_451_io_o_g;
  wire  Black_451_io_o_p;
  Black Black_451 (
    .io_i_pj(Black_451_io_i_pj),
    .io_i_gj(Black_451_io_i_gj),
    .io_i_pk(Black_451_io_i_pk),
    .io_i_gk(Black_451_io_i_gk),
    .io_o_g(Black_451_io_o_g),
    .io_o_p(Black_451_io_o_p)
  );

  wire  Black_458_io_i_pj;
  wire  Black_458_io_i_gj;
  wire  Black_458_io_i_pk;
  wire  Black_458_io_i_gk;
  wire  Black_458_io_o_g;
  wire  Black_458_io_o_p;
  Black Black_458 (
    .io_i_pj(Black_458_io_i_pj),
    .io_i_gj(Black_458_io_i_gj),
    .io_i_pk(Black_458_io_i_pk),
    .io_i_gk(Black_458_io_i_gk),
    .io_o_g(Black_458_io_o_g),
    .io_o_p(Black_458_io_o_p)
  );

  wire  Black_461_io_i_pj;
  wire  Black_461_io_i_gj;
  wire  Black_461_io_i_pk;
  wire  Black_461_io_i_gk;
  wire  Black_461_io_o_g;
  wire  Black_461_io_o_p;
  Black Black_461 (
    .io_i_pj(Black_461_io_i_pj),
    .io_i_gj(Black_461_io_i_gj),
    .io_i_pk(Black_461_io_i_pk),
    .io_i_gk(Black_461_io_i_gk),
    .io_o_g(Black_461_io_o_g),
    .io_o_p(Black_461_io_o_p)
  );

  wire  PG_462_io_i_a;
  wire  PG_462_io_i_b;
  wire  PG_462_io_o_p;
  wire  PG_462_io_o_g;
  PG PG_462 (
    .io_i_a(PG_462_io_i_a),
    .io_i_b(PG_462_io_i_b),
    .io_o_p(PG_462_io_o_p),
    .io_o_g(PG_462_io_o_g)
  );

  wire  Black_463_io_i_pj;
  wire  Black_463_io_i_gj;
  wire  Black_463_io_i_pk;
  wire  Black_463_io_i_gk;
  wire  Black_463_io_o_g;
  wire  Black_463_io_o_p;
  Black Black_463 (
    .io_i_pj(Black_463_io_i_pj),
    .io_i_gj(Black_463_io_i_gj),
    .io_i_pk(Black_463_io_i_pk),
    .io_i_gk(Black_463_io_i_gk),
    .io_o_g(Black_463_io_o_g),
    .io_o_p(Black_463_io_o_p)
  );

  wire  Black_464_io_i_pj;
  wire  Black_464_io_i_gj;
  wire  Black_464_io_i_pk;
  wire  Black_464_io_i_gk;
  wire  Black_464_io_o_g;
  wire  Black_464_io_o_p;
  Black Black_464 (
    .io_i_pj(Black_464_io_i_pj),
    .io_i_gj(Black_464_io_i_gj),
    .io_i_pk(Black_464_io_i_pk),
    .io_i_gk(Black_464_io_i_gk),
    .io_o_g(Black_464_io_o_g),
    .io_o_p(Black_464_io_o_p)
  );

  wire  Black_467_io_i_pj;
  wire  Black_467_io_i_gj;
  wire  Black_467_io_i_pk;
  wire  Black_467_io_i_gk;
  wire  Black_467_io_o_g;
  wire  Black_467_io_o_p;
  Black Black_467 (
    .io_i_pj(Black_467_io_i_pj),
    .io_i_gj(Black_467_io_i_gj),
    .io_i_pk(Black_467_io_i_pk),
    .io_i_gk(Black_467_io_i_gk),
    .io_o_g(Black_467_io_o_g),
    .io_o_p(Black_467_io_o_p)
  );

  wire  Black_469_io_i_pj;
  wire  Black_469_io_i_gj;
  wire  Black_469_io_i_pk;
  wire  Black_469_io_i_gk;
  wire  Black_469_io_o_g;
  wire  Black_469_io_o_p;
  Black Black_469 (
    .io_i_pj(Black_469_io_i_pj),
    .io_i_gj(Black_469_io_i_gj),
    .io_i_pk(Black_469_io_i_pk),
    .io_i_gk(Black_469_io_i_gk),
    .io_o_g(Black_469_io_o_g),
    .io_o_p(Black_469_io_o_p)
  );

  wire  Black_472_io_i_pj;
  wire  Black_472_io_i_gj;
  wire  Black_472_io_i_pk;
  wire  Black_472_io_i_gk;
  wire  Black_472_io_o_g;
  wire  Black_472_io_o_p;
  Black Black_472 (
    .io_i_pj(Black_472_io_i_pj),
    .io_i_gj(Black_472_io_i_gj),
    .io_i_pk(Black_472_io_i_pk),
    .io_i_gk(Black_472_io_i_gk),
    .io_o_g(Black_472_io_o_g),
    .io_o_p(Black_472_io_o_p)
  );

  wire  PG_473_io_i_a;
  wire  PG_473_io_i_b;
  wire  PG_473_io_o_p;
  wire  PG_473_io_o_g;
  PG PG_473 (
    .io_i_a(PG_473_io_i_a),
    .io_i_b(PG_473_io_i_b),
    .io_o_p(PG_473_io_o_p),
    .io_o_g(PG_473_io_o_g)
  );

  wire  Black_478_io_i_pj;
  wire  Black_478_io_i_gj;
  wire  Black_478_io_i_pk;
  wire  Black_478_io_i_gk;
  wire  Black_478_io_o_g;
  wire  Black_478_io_o_p;
  Black Black_478 (
    .io_i_pj(Black_478_io_i_pj),
    .io_i_gj(Black_478_io_i_gj),
    .io_i_pk(Black_478_io_i_pk),
    .io_i_gk(Black_478_io_i_gk),
    .io_o_g(Black_478_io_o_g),
    .io_o_p(Black_478_io_o_p)
  );

  wire  Black_479_io_i_pj;
  wire  Black_479_io_i_gj;
  wire  Black_479_io_i_pk;
  wire  Black_479_io_i_gk;
  wire  Black_479_io_o_g;
  wire  Black_479_io_o_p;
  Black Black_479 (
    .io_i_pj(Black_479_io_i_pj),
    .io_i_gj(Black_479_io_i_gj),
    .io_i_pk(Black_479_io_i_pk),
    .io_i_gk(Black_479_io_i_gk),
    .io_o_g(Black_479_io_o_g),
    .io_o_p(Black_479_io_o_p)
  );

  wire  Black_482_io_i_pj;
  wire  Black_482_io_i_gj;
  wire  Black_482_io_i_pk;
  wire  Black_482_io_i_gk;
  wire  Black_482_io_o_g;
  wire  Black_482_io_o_p;
  Black Black_482 (
    .io_i_pj(Black_482_io_i_pj),
    .io_i_gj(Black_482_io_i_gj),
    .io_i_pk(Black_482_io_i_pk),
    .io_i_gk(Black_482_io_i_gk),
    .io_o_g(Black_482_io_o_g),
    .io_o_p(Black_482_io_o_p)
  );

  wire  PG_483_io_i_a;
  wire  PG_483_io_i_b;
  wire  PG_483_io_o_p;
  wire  PG_483_io_o_g;
  PG PG_483 (
    .io_i_a(PG_483_io_i_a),
    .io_i_b(PG_483_io_i_b),
    .io_o_p(PG_483_io_o_p),
    .io_o_g(PG_483_io_o_g)
  );

  wire  Black_486_io_i_pj;
  wire  Black_486_io_i_gj;
  wire  Black_486_io_i_pk;
  wire  Black_486_io_i_gk;
  wire  Black_486_io_o_g;
  wire  Black_486_io_o_p;
  Black Black_486 (
    .io_i_pj(Black_486_io_i_pj),
    .io_i_gj(Black_486_io_i_gj),
    .io_i_pk(Black_486_io_i_pk),
    .io_i_gk(Black_486_io_i_gk),
    .io_o_g(Black_486_io_o_g),
    .io_o_p(Black_486_io_o_p)
  );

  wire  Black_487_io_i_pj;
  wire  Black_487_io_i_gj;
  wire  Black_487_io_i_pk;
  wire  Black_487_io_i_gk;
  wire  Black_487_io_o_g;
  wire  Black_487_io_o_p;
  Black Black_487 (
    .io_i_pj(Black_487_io_i_pj),
    .io_i_gj(Black_487_io_i_gj),
    .io_i_pk(Black_487_io_i_pk),
    .io_i_gk(Black_487_io_i_gk),
    .io_o_g(Black_487_io_o_g),
    .io_o_p(Black_487_io_o_p)
  );

  wire  Black_491_io_i_pj;
  wire  Black_491_io_i_gj;
  wire  Black_491_io_i_pk;
  wire  Black_491_io_i_gk;
  wire  Black_491_io_o_g;
  wire  Black_491_io_o_p;
  Black Black_491 (
    .io_i_pj(Black_491_io_i_pj),
    .io_i_gj(Black_491_io_i_gj),
    .io_i_pk(Black_491_io_i_pk),
    .io_i_gk(Black_491_io_i_gk),
    .io_o_g(Black_491_io_o_g),
    .io_o_p(Black_491_io_o_p)
  );

  wire  PG_492_io_i_a;
  wire  PG_492_io_i_b;
  wire  PG_492_io_o_p;
  wire  PG_492_io_o_g;
  PG PG_492 (
    .io_i_a(PG_492_io_i_a),
    .io_i_b(PG_492_io_i_b),
    .io_o_p(PG_492_io_o_p),
    .io_o_g(PG_492_io_o_g)
  );

  wire  Black_493_io_i_pj;
  wire  Black_493_io_i_gj;
  wire  Black_493_io_i_pk;
  wire  Black_493_io_i_gk;
  wire  Black_493_io_o_g;
  wire  Black_493_io_o_p;
  Black Black_493 (
    .io_i_pj(Black_493_io_i_pj),
    .io_i_gj(Black_493_io_i_gj),
    .io_i_pk(Black_493_io_i_pk),
    .io_i_gk(Black_493_io_i_gk),
    .io_o_g(Black_493_io_o_g),
    .io_o_p(Black_493_io_o_p)
  );

  wire  Black_494_io_i_pj;
  wire  Black_494_io_i_gj;
  wire  Black_494_io_i_pk;
  wire  Black_494_io_i_gk;
  wire  Black_494_io_o_g;
  wire  Black_494_io_o_p;
  Black Black_494 (
    .io_i_pj(Black_494_io_i_pj),
    .io_i_gj(Black_494_io_i_gj),
    .io_i_pk(Black_494_io_i_pk),
    .io_i_gk(Black_494_io_i_gk),
    .io_o_g(Black_494_io_o_g),
    .io_o_p(Black_494_io_o_p)
  );

  wire  Black_495_io_i_pj;
  wire  Black_495_io_i_gj;
  wire  Black_495_io_i_pk;
  wire  Black_495_io_i_gk;
  wire  Black_495_io_o_g;
  wire  Black_495_io_o_p;
  Black Black_495 (
    .io_i_pj(Black_495_io_i_pj),
    .io_i_gj(Black_495_io_i_gj),
    .io_i_pk(Black_495_io_i_pk),
    .io_i_gk(Black_495_io_i_gk),
    .io_o_g(Black_495_io_o_g),
    .io_o_p(Black_495_io_o_p)
  );

  wire  Black_497_io_i_pj;
  wire  Black_497_io_i_gj;
  wire  Black_497_io_i_pk;
  wire  Black_497_io_i_gk;
  wire  Black_497_io_o_g;
  wire  Black_497_io_o_p;
  Black Black_497 (
    .io_i_pj(Black_497_io_i_pj),
    .io_i_gj(Black_497_io_i_gj),
    .io_i_pk(Black_497_io_i_pk),
    .io_i_gk(Black_497_io_i_gk),
    .io_o_g(Black_497_io_o_g),
    .io_o_p(Black_497_io_o_p)
  );

  wire  Black_498_io_i_pj;
  wire  Black_498_io_i_gj;
  wire  Black_498_io_i_pk;
  wire  Black_498_io_i_gk;
  wire  Black_498_io_o_g;
  wire  Black_498_io_o_p;
  Black Black_498 (
    .io_i_pj(Black_498_io_i_pj),
    .io_i_gj(Black_498_io_i_gj),
    .io_i_pk(Black_498_io_i_pk),
    .io_i_gk(Black_498_io_i_gk),
    .io_o_g(Black_498_io_o_g),
    .io_o_p(Black_498_io_o_p)
  );

  wire  Black_499_io_i_pj;
  wire  Black_499_io_i_gj;
  wire  Black_499_io_i_pk;
  wire  Black_499_io_i_gk;
  wire  Black_499_io_o_g;
  wire  Black_499_io_o_p;
  Black Black_499 (
    .io_i_pj(Black_499_io_i_pj),
    .io_i_gj(Black_499_io_i_gj),
    .io_i_pk(Black_499_io_i_pk),
    .io_i_gk(Black_499_io_i_gk),
    .io_o_g(Black_499_io_o_g),
    .io_o_p(Black_499_io_o_p)
  );

  wire  PG_500_io_i_a;
  wire  PG_500_io_i_b;
  wire  PG_500_io_o_p;
  wire  PG_500_io_o_g;
  PG PG_500 (
    .io_i_a(PG_500_io_i_a),
    .io_i_b(PG_500_io_i_b),
    .io_o_p(PG_500_io_o_p),
    .io_o_g(PG_500_io_o_g)
  );

  wire  Black_502_io_i_pj;
  wire  Black_502_io_i_gj;
  wire  Black_502_io_i_pk;
  wire  Black_502_io_i_gk;
  wire  Black_502_io_o_g;
  wire  Black_502_io_o_p;
  Black Black_502 (
    .io_i_pj(Black_502_io_i_pj),
    .io_i_gj(Black_502_io_i_gj),
    .io_i_pk(Black_502_io_i_pk),
    .io_i_gk(Black_502_io_i_gk),
    .io_o_g(Black_502_io_o_g),
    .io_o_p(Black_502_io_o_p)
  );

  wire  Black_503_io_i_pj;
  wire  Black_503_io_i_gj;
  wire  Black_503_io_i_pk;
  wire  Black_503_io_i_gk;
  wire  Black_503_io_o_g;
  wire  Black_503_io_o_p;
  Black Black_503 (
    .io_i_pj(Black_503_io_i_pj),
    .io_i_gj(Black_503_io_i_gj),
    .io_i_pk(Black_503_io_i_pk),
    .io_i_gk(Black_503_io_i_gk),
    .io_o_g(Black_503_io_o_g),
    .io_o_p(Black_503_io_o_p)
  );

  wire  Black_506_io_i_pj;
  wire  Black_506_io_i_gj;
  wire  Black_506_io_i_pk;
  wire  Black_506_io_i_gk;
  wire  Black_506_io_o_g;
  wire  Black_506_io_o_p;
  Black Black_506 (
    .io_i_pj(Black_506_io_i_pj),
    .io_i_gj(Black_506_io_i_gj),
    .io_i_pk(Black_506_io_i_pk),
    .io_i_gk(Black_506_io_i_gk),
    .io_o_g(Black_506_io_o_g),
    .io_o_p(Black_506_io_o_p)
  );

  wire  PG_507_io_i_a;
  wire  PG_507_io_i_b;
  wire  PG_507_io_o_p;
  wire  PG_507_io_o_g;
  PG PG_507 (
    .io_i_a(PG_507_io_i_a),
    .io_i_b(PG_507_io_i_b),
    .io_o_p(PG_507_io_o_p),
    .io_o_g(PG_507_io_o_g)
  );

  wire  Black_508_io_i_pj;
  wire  Black_508_io_i_gj;
  wire  Black_508_io_i_pk;
  wire  Black_508_io_i_gk;
  wire  Black_508_io_o_g;
  wire  Black_508_io_o_p;
  Black Black_508 (
    .io_i_pj(Black_508_io_i_pj),
    .io_i_gj(Black_508_io_i_gj),
    .io_i_pk(Black_508_io_i_pk),
    .io_i_gk(Black_508_io_i_gk),
    .io_o_g(Black_508_io_o_g),
    .io_o_p(Black_508_io_o_p)
  );

  wire  Black_512_io_i_pj;
  wire  Black_512_io_i_gj;
  wire  Black_512_io_i_pk;
  wire  Black_512_io_i_gk;
  wire  Black_512_io_o_g;
  wire  Black_512_io_o_p;
  Black Black_512 (
    .io_i_pj(Black_512_io_i_pj),
    .io_i_gj(Black_512_io_i_gj),
    .io_i_pk(Black_512_io_i_pk),
    .io_i_gk(Black_512_io_i_gk),
    .io_o_g(Black_512_io_o_g),
    .io_o_p(Black_512_io_o_p)
  );

  wire  PG_513_io_i_a;
  wire  PG_513_io_i_b;
  wire  PG_513_io_o_p;
  wire  PG_513_io_o_g;
  PG PG_513 (
    .io_i_a(PG_513_io_i_a),
    .io_i_b(PG_513_io_i_b),
    .io_o_p(PG_513_io_o_p),
    .io_o_g(PG_513_io_o_g)
  );

  wire  Black_514_io_i_pj;
  wire  Black_514_io_i_gj;
  wire  Black_514_io_i_pk;
  wire  Black_514_io_i_gk;
  wire  Black_514_io_o_g;
  wire  Black_514_io_o_p;
  Black Black_514 (
    .io_i_pj(Black_514_io_i_pj),
    .io_i_gj(Black_514_io_i_gj),
    .io_i_pk(Black_514_io_i_pk),
    .io_i_gk(Black_514_io_i_gk),
    .io_o_g(Black_514_io_o_g),
    .io_o_p(Black_514_io_o_p)
  );

  wire  Black_515_io_i_pj;
  wire  Black_515_io_i_gj;
  wire  Black_515_io_i_pk;
  wire  Black_515_io_i_gk;
  wire  Black_515_io_o_g;
  wire  Black_515_io_o_p;
  Black Black_515 (
    .io_i_pj(Black_515_io_i_pj),
    .io_i_gj(Black_515_io_i_gj),
    .io_i_pk(Black_515_io_i_pk),
    .io_i_gk(Black_515_io_i_gk),
    .io_o_g(Black_515_io_o_g),
    .io_o_p(Black_515_io_o_p)
  );

  wire  Black_517_io_i_pj;
  wire  Black_517_io_i_gj;
  wire  Black_517_io_i_pk;
  wire  Black_517_io_i_gk;
  wire  Black_517_io_o_g;
  wire  Black_517_io_o_p;
  Black Black_517 (
    .io_i_pj(Black_517_io_i_pj),
    .io_i_gj(Black_517_io_i_gj),
    .io_i_pk(Black_517_io_i_pk),
    .io_i_gk(Black_517_io_i_gk),
    .io_o_g(Black_517_io_o_g),
    .io_o_p(Black_517_io_o_p)
  );

  wire  PG_518_io_i_a;
  wire  PG_518_io_i_b;
  wire  PG_518_io_o_p;
  wire  PG_518_io_o_g;
  PG PG_518 (
    .io_i_a(PG_518_io_i_a),
    .io_i_b(PG_518_io_i_b),
    .io_o_p(PG_518_io_o_p),
    .io_o_g(PG_518_io_o_g)
  );

  wire  Black_519_io_i_pj;
  wire  Black_519_io_i_gj;
  wire  Black_519_io_i_pk;
  wire  Black_519_io_i_gk;
  wire  Black_519_io_o_g;
  wire  Black_519_io_o_p;
  Black Black_519 (
    .io_i_pj(Black_519_io_i_pj),
    .io_i_gj(Black_519_io_i_gj),
    .io_i_pk(Black_519_io_i_pk),
    .io_i_gk(Black_519_io_i_gk),
    .io_o_g(Black_519_io_o_g),
    .io_o_p(Black_519_io_o_p)
  );

  wire  Black_521_io_i_pj;
  wire  Black_521_io_i_gj;
  wire  Black_521_io_i_pk;
  wire  Black_521_io_i_gk;
  wire  Black_521_io_o_g;
  wire  Black_521_io_o_p;
  Black Black_521 (
    .io_i_pj(Black_521_io_i_pj),
    .io_i_gj(Black_521_io_i_gj),
    .io_i_pk(Black_521_io_i_pk),
    .io_i_gk(Black_521_io_i_gk),
    .io_o_g(Black_521_io_o_g),
    .io_o_p(Black_521_io_o_p)
  );

  wire  PG_522_io_i_a;
  wire  PG_522_io_i_b;
  wire  PG_522_io_o_p;
  wire  PG_522_io_o_g;
  PG PG_522 (
    .io_i_a(PG_522_io_i_a),
    .io_i_b(PG_522_io_i_b),
    .io_o_p(PG_522_io_o_p),
    .io_o_g(PG_522_io_o_g)
  );

  wire  Black_523_io_i_pj;
  wire  Black_523_io_i_gj;
  wire  Black_523_io_i_pk;
  wire  Black_523_io_i_gk;
  wire  Black_523_io_o_g;
  wire  Black_523_io_o_p;
  Black Black_523 (
    .io_i_pj(Black_523_io_i_pj),
    .io_i_gj(Black_523_io_i_gj),
    .io_i_pk(Black_523_io_i_pk),
    .io_i_gk(Black_523_io_i_gk),
    .io_o_g(Black_523_io_o_g),
    .io_o_p(Black_523_io_o_p)
  );

  wire  Black_524_io_i_pj;
  wire  Black_524_io_i_gj;
  wire  Black_524_io_i_pk;
  wire  Black_524_io_i_gk;
  wire  Black_524_io_o_g;
  wire  Black_524_io_o_p;
  Black Black_524 (
    .io_i_pj(Black_524_io_i_pj),
    .io_i_gj(Black_524_io_i_gj),
    .io_i_pk(Black_524_io_i_pk),
    .io_i_gk(Black_524_io_i_gk),
    .io_o_g(Black_524_io_o_g),
    .io_o_p(Black_524_io_o_p)
  );

  wire  PG_525_io_i_a;
  wire  PG_525_io_i_b;
  wire  PG_525_io_o_p;
  wire  PG_525_io_o_g;
  PG PG_525 (
    .io_i_a(PG_525_io_i_a),
    .io_i_b(PG_525_io_i_b),
    .io_o_p(PG_525_io_o_p),
    .io_o_g(PG_525_io_o_g)
  );

  wire  Black_526_io_i_pj;
  wire  Black_526_io_i_gj;
  wire  Black_526_io_i_pk;
  wire  Black_526_io_i_gk;
  wire  Black_526_io_o_g;
  wire  Black_526_io_o_p;
  Black Black_526 (
    .io_i_pj(Black_526_io_i_pj),
    .io_i_gj(Black_526_io_i_gj),
    .io_i_pk(Black_526_io_i_pk),
    .io_i_gk(Black_526_io_i_gk),
    .io_o_g(Black_526_io_o_g),
    .io_o_p(Black_526_io_o_p)
  );

  wire  PG_527_io_i_a;
  wire  PG_527_io_i_b;
  wire  PG_527_io_o_p;
  wire  PG_527_io_o_g;
  PG PG_527 (
    .io_i_a(PG_527_io_i_a),
    .io_i_b(PG_527_io_i_b),
    .io_o_p(PG_527_io_o_p),
    .io_o_g(PG_527_io_o_g)
  );

  wire  res_0 = PG_527_io_o_p;

  wire  res_1 = PG_525_io_o_p ^ PG_527_io_o_g;

  wire  res_2 = PG_522_io_o_p ^ Black_526_io_o_g;

  wire  res_3 = PG_518_io_o_p ^ Black_524_io_o_g;

  wire  res_4 = PG_513_io_o_p ^ Black_521_io_o_g;

  wire  res_5 = PG_507_io_o_p ^ Black_517_io_o_g;

  wire  res_6 = PG_500_io_o_p ^ Black_512_io_o_g;

  wire  res_7 = PG_492_io_o_p ^ Black_506_io_o_g;

  wire  res_8 = PG_483_io_o_p ^ Black_499_io_o_g;

  wire  res_9 = PG_473_io_o_p ^ Black_491_io_o_g;

  wire  res_10 = PG_462_io_o_p ^ Black_482_io_o_g;

  wire  res_11 = PG_450_io_o_p ^ Black_472_io_o_g;

  wire  res_12 = PG_437_io_o_p ^ Black_461_io_o_g;

  wire  res_13 = PG_423_io_o_p ^ Black_449_io_o_g;

  wire  res_14 = PG_408_io_o_p ^ Black_436_io_o_g;

  wire  res_15 = PG_392_io_o_p ^ Black_422_io_o_g;

  wire  res_16 = PG_375_io_o_p ^ Black_407_io_o_g;

  wire  res_17 = PG_357_io_o_p ^ Black_391_io_o_g;

  wire  res_18 = PG_338_io_o_p ^ Black_374_io_o_g;

  wire  res_19 = PG_318_io_o_p ^ Black_356_io_o_g;

  wire  res_20 = PG_297_io_o_p ^ Black_337_io_o_g;

  wire  res_21 = PG_275_io_o_p ^ Black_317_io_o_g;

  wire  res_22 = PG_252_io_o_p ^ Black_296_io_o_g;

  wire  res_23 = PG_228_io_o_p ^ Black_274_io_o_g;

  wire  res_24 = PG_203_io_o_p ^ Black_251_io_o_g;

  wire  res_25 = PG_177_io_o_p ^ Black_227_io_o_g;

  wire  res_26 = PG_150_io_o_p ^ Black_202_io_o_g;

  wire  res_27 = PG_122_io_o_p ^ Black_176_io_o_g;

  wire  res_28 = PG_93_io_o_p ^ Black_149_io_o_g;

  wire  res_29 = PG_63_io_o_p ^ Black_121_io_o_g;

  wire  res_30 = PG_32_io_o_p ^ Black_92_io_o_g;

  wire  res_31 = PG_0_io_o_p ^ Black_62_io_o_g;
assign io_outs = {res_31, res_30, res_29, res_28, res_27, res_26, res_25, res_24, res_23, res_22, res_21, res_20, res_19, res_18, res_17, res_16, res_15, res_14, res_13, res_12, res_11, res_10, res_9, res_8, res_7, res_6, res_5, res_4, res_3, res_2, res_1, res_0};

  assign PG_527_io_i_a = io_augend[0];
  assign PG_527_io_i_b = io_addend[0];

  assign PG_525_io_i_a = io_augend[1];
  assign PG_525_io_i_b = io_addend[1];

  assign PG_522_io_i_a = io_augend[2];
  assign PG_522_io_i_b = io_addend[2];

  assign PG_518_io_i_a = io_augend[3];
  assign PG_518_io_i_b = io_addend[3];

  assign PG_513_io_i_a = io_augend[4];
  assign PG_513_io_i_b = io_addend[4];

  assign PG_507_io_i_a = io_augend[5];
  assign PG_507_io_i_b = io_addend[5];

  assign PG_500_io_i_a = io_augend[6];
  assign PG_500_io_i_b = io_addend[6];

  assign PG_492_io_i_a = io_augend[7];
  assign PG_492_io_i_b = io_addend[7];

  assign PG_483_io_i_a = io_augend[8];
  assign PG_483_io_i_b = io_addend[8];

  assign PG_473_io_i_a = io_augend[9];
  assign PG_473_io_i_b = io_addend[9];

  assign PG_462_io_i_a = io_augend[10];
  assign PG_462_io_i_b = io_addend[10];

  assign PG_450_io_i_a = io_augend[11];
  assign PG_450_io_i_b = io_addend[11];

  assign PG_437_io_i_a = io_augend[12];
  assign PG_437_io_i_b = io_addend[12];

  assign PG_423_io_i_a = io_augend[13];
  assign PG_423_io_i_b = io_addend[13];

  assign PG_408_io_i_a = io_augend[14];
  assign PG_408_io_i_b = io_addend[14];

  assign PG_392_io_i_a = io_augend[15];
  assign PG_392_io_i_b = io_addend[15];

  assign PG_375_io_i_a = io_augend[16];
  assign PG_375_io_i_b = io_addend[16];

  assign PG_357_io_i_a = io_augend[17];
  assign PG_357_io_i_b = io_addend[17];

  assign PG_338_io_i_a = io_augend[18];
  assign PG_338_io_i_b = io_addend[18];

  assign PG_318_io_i_a = io_augend[19];
  assign PG_318_io_i_b = io_addend[19];

  assign PG_297_io_i_a = io_augend[20];
  assign PG_297_io_i_b = io_addend[20];

  assign PG_275_io_i_a = io_augend[21];
  assign PG_275_io_i_b = io_addend[21];

  assign PG_252_io_i_a = io_augend[22];
  assign PG_252_io_i_b = io_addend[22];

  assign PG_228_io_i_a = io_augend[23];
  assign PG_228_io_i_b = io_addend[23];

  assign PG_203_io_i_a = io_augend[24];
  assign PG_203_io_i_b = io_addend[24];

  assign PG_177_io_i_a = io_augend[25];
  assign PG_177_io_i_b = io_addend[25];

  assign PG_150_io_i_a = io_augend[26];
  assign PG_150_io_i_b = io_addend[26];

  assign PG_122_io_i_a = io_augend[27];
  assign PG_122_io_i_b = io_addend[27];

  assign PG_93_io_i_a = io_augend[28];
  assign PG_93_io_i_b = io_addend[28];

  assign PG_63_io_i_a = io_augend[29];
  assign PG_63_io_i_b = io_addend[29];

  assign PG_32_io_i_a = io_augend[30];
  assign PG_32_io_i_b = io_addend[30];

  assign PG_0_io_i_a = io_augend[31];
  assign PG_0_io_i_b = io_addend[31];

  assign Black_1_io_i_pj = PG_32_io_o_p;
  assign Black_1_io_i_gj = PG_32_io_o_g;
  assign Black_1_io_i_pk = PG_0_io_o_p;
  assign Black_1_io_i_gk = PG_0_io_o_g;

  assign Black_3_io_i_pj = Black_64_io_o_p;
  assign Black_3_io_i_gj = Black_64_io_o_g;
  assign Black_3_io_i_pk = Black_1_io_o_p;
  assign Black_3_io_i_gk = Black_1_io_o_g;

  assign Black_7_io_i_pj = Black_125_io_o_p;
  assign Black_7_io_i_gj = Black_125_io_o_g;
  assign Black_7_io_i_pk = Black_3_io_o_p;
  assign Black_7_io_i_gk = Black_3_io_o_g;

  assign Black_15_io_i_pj = Black_235_io_o_p;
  assign Black_15_io_i_gj = Black_235_io_o_g;
  assign Black_15_io_i_pk = Black_7_io_o_p;
  assign Black_15_io_i_gk = Black_7_io_o_g;

  assign Black_31_io_i_pj = Black_407_io_o_p;
  assign Black_31_io_i_gj = Black_407_io_o_g;
  assign Black_31_io_i_pk = Black_15_io_o_p;
  assign Black_31_io_i_gk = Black_15_io_o_g;

  assign Black_34_io_i_pj = Black_64_io_o_p;
  assign Black_34_io_i_gj = Black_64_io_o_g;
  assign Black_34_io_i_pk = PG_32_io_o_p;
  assign Black_34_io_i_gk = PG_32_io_o_g;

  assign Black_38_io_i_pj = Black_125_io_o_p;
  assign Black_38_io_i_gj = Black_125_io_o_g;
  assign Black_38_io_i_pk = Black_34_io_o_p;
  assign Black_38_io_i_gk = Black_34_io_o_g;

  assign Black_46_io_i_pj = Black_235_io_o_p;
  assign Black_46_io_i_gj = Black_235_io_o_g;
  assign Black_46_io_i_pk = Black_38_io_o_p;
  assign Black_46_io_i_gk = Black_38_io_o_g;

  assign Black_53_io_i_pj = Black_398_io_o_p;
  assign Black_53_io_i_gj = Black_398_io_o_g;
  assign Black_53_io_i_pk = Black_46_io_o_p;
  assign Black_53_io_i_gk = Black_46_io_o_g;

  assign Black_62_io_i_pj = Black_491_io_o_p;
  assign Black_62_io_i_gj = Black_491_io_o_g;
  assign Black_62_io_i_pk = Black_53_io_o_p;
  assign Black_62_io_i_gk = Black_53_io_o_g;

  assign Black_64_io_i_pj = PG_93_io_o_p;
  assign Black_64_io_i_gj = PG_93_io_o_g;
  assign Black_64_io_i_pk = PG_63_io_o_p;
  assign Black_64_io_i_gk = PG_63_io_o_g;

  assign Black_68_io_i_pj = Black_125_io_o_p;
  assign Black_68_io_i_gj = Black_125_io_o_g;
  assign Black_68_io_i_pk = Black_64_io_o_p;
  assign Black_68_io_i_gk = Black_64_io_o_g;

  assign Black_87_io_i_pj = Black_246_io_o_p;
  assign Black_87_io_i_gj = Black_246_io_o_g;
  assign Black_87_io_i_pk = Black_68_io_o_p;
  assign Black_87_io_i_gk = Black_68_io_o_g;

  assign Black_90_io_i_pj = Black_515_io_o_p;
  assign Black_90_io_i_gj = Black_515_io_o_g;
  assign Black_90_io_i_pk = Black_87_io_o_p;
  assign Black_90_io_i_gk = Black_87_io_o_g;

  assign Black_92_io_i_pj = Black_526_io_o_p;
  assign Black_92_io_i_gj = Black_526_io_o_g;
  assign Black_92_io_i_pk = Black_90_io_o_p;
  assign Black_92_io_i_gk = Black_90_io_o_g;

  assign Black_99_io_i_pj = Black_127_io_o_p;
  assign Black_99_io_i_gj = Black_127_io_o_g;
  assign Black_99_io_i_pk = PG_93_io_o_p;
  assign Black_99_io_i_gk = PG_93_io_o_g;

  assign Black_105_io_i_pj = Black_280_io_o_p;
  assign Black_105_io_i_gj = Black_280_io_o_g;
  assign Black_105_io_i_pk = Black_99_io_o_p;
  assign Black_105_io_i_gk = Black_99_io_o_g;

  assign Black_121_io_i_pj = Black_407_io_o_p;
  assign Black_121_io_i_gj = Black_407_io_o_g;
  assign Black_121_io_i_pk = Black_105_io_o_p;
  assign Black_121_io_i_gk = Black_105_io_o_g;

  assign Black_123_io_i_pj = PG_150_io_o_p;
  assign Black_123_io_i_gj = PG_150_io_o_g;
  assign Black_123_io_i_pk = PG_122_io_o_p;
  assign Black_123_io_i_gk = PG_122_io_o_g;

  assign Black_125_io_i_pj = Black_178_io_o_p;
  assign Black_125_io_i_gj = Black_178_io_o_g;
  assign Black_125_io_i_pk = Black_123_io_o_p;
  assign Black_125_io_i_gk = Black_123_io_o_g;

  assign Black_127_io_i_pj = Black_229_io_o_p;
  assign Black_127_io_i_gj = Black_229_io_o_g;
  assign Black_127_io_i_pk = Black_125_io_o_p;
  assign Black_127_io_i_gk = Black_125_io_o_g;

  assign Black_133_io_i_pj = Black_280_io_o_p;
  assign Black_133_io_i_gj = Black_280_io_o_g;
  assign Black_133_io_i_pk = Black_127_io_o_p;
  assign Black_133_io_i_gk = Black_127_io_o_g;

  assign Black_135_io_i_pj = Black_393_io_o_p;
  assign Black_135_io_i_gj = Black_393_io_o_g;
  assign Black_135_io_i_pk = Black_133_io_o_p;
  assign Black_135_io_i_gk = Black_133_io_o_g;

  assign Black_145_io_i_pj = Black_432_io_o_p;
  assign Black_145_io_i_gj = Black_432_io_o_g;
  assign Black_145_io_i_pk = Black_135_io_o_p;
  assign Black_145_io_i_gk = Black_135_io_o_g;

  assign Black_149_io_i_pj = Black_521_io_o_p;
  assign Black_149_io_i_gj = Black_521_io_o_g;
  assign Black_149_io_i_pk = Black_145_io_o_p;
  assign Black_149_io_i_gk = Black_145_io_o_g;

  assign Black_152_io_i_pj = Black_178_io_o_p;
  assign Black_152_io_i_gj = Black_178_io_o_g;
  assign Black_152_io_i_pk = PG_150_io_o_p;
  assign Black_152_io_i_gk = PG_150_io_o_g;

  assign Black_153_io_i_pj = PG_228_io_o_p;
  assign Black_153_io_i_gj = PG_228_io_o_g;
  assign Black_153_io_i_pk = Black_152_io_o_p;
  assign Black_153_io_i_gk = Black_152_io_o_g;

  assign Black_160_io_i_pj = Black_258_io_o_p;
  assign Black_160_io_i_gj = Black_258_io_o_g;
  assign Black_160_io_i_pk = Black_153_io_o_p;
  assign Black_160_io_i_gk = Black_153_io_o_g;

  assign Black_162_io_i_pj = Black_393_io_o_p;
  assign Black_162_io_i_gj = Black_393_io_o_g;
  assign Black_162_io_i_pk = Black_160_io_o_p;
  assign Black_162_io_i_gk = Black_160_io_o_g;

  assign Black_176_io_i_pj = Black_436_io_o_p;
  assign Black_176_io_i_gj = Black_436_io_o_g;
  assign Black_176_io_i_pk = Black_162_io_o_p;
  assign Black_176_io_i_gk = Black_162_io_o_g;

  assign Black_178_io_i_pj = PG_203_io_o_p;
  assign Black_178_io_i_gj = PG_203_io_o_g;
  assign Black_178_io_i_pk = PG_177_io_o_p;
  assign Black_178_io_i_gk = PG_177_io_o_g;

  assign Black_180_io_i_pj = Black_229_io_o_p;
  assign Black_180_io_i_gj = Black_229_io_o_g;
  assign Black_180_io_i_pk = Black_178_io_o_p;
  assign Black_180_io_i_gk = Black_178_io_o_g;

  assign Black_202_io_i_pj = Black_296_io_o_p;
  assign Black_202_io_i_gj = Black_296_io_o_g;
  assign Black_202_io_i_pk = Black_180_io_o_p;
  assign Black_202_io_i_gk = Black_180_io_o_g;

  assign Black_211_io_i_pj = Black_235_io_o_p;
  assign Black_211_io_i_gj = Black_235_io_o_g;
  assign Black_211_io_i_pk = PG_203_io_o_p;
  assign Black_211_io_i_gk = PG_203_io_o_g;

  assign Black_227_io_i_pj = Black_407_io_o_p;
  assign Black_227_io_i_gj = Black_407_io_o_g;
  assign Black_227_io_i_pk = Black_211_io_o_p;
  assign Black_227_io_i_gk = Black_211_io_o_g;

  assign Black_229_io_i_pj = PG_252_io_o_p;
  assign Black_229_io_i_gj = PG_252_io_o_g;
  assign Black_229_io_i_pk = PG_228_io_o_p;
  assign Black_229_io_i_gk = PG_228_io_o_g;

  assign Black_231_io_i_pj = Black_276_io_o_p;
  assign Black_231_io_i_gj = Black_276_io_o_g;
  assign Black_231_io_i_pk = Black_229_io_o_p;
  assign Black_231_io_i_gk = Black_229_io_o_g;

  assign Black_235_io_i_pj = Black_321_io_o_p;
  assign Black_235_io_i_gj = Black_321_io_o_g;
  assign Black_235_io_i_pk = Black_231_io_o_p;
  assign Black_235_io_i_gk = Black_231_io_o_g;

  assign Black_238_io_i_pj = Black_394_io_o_p;
  assign Black_238_io_i_gj = Black_394_io_o_g;
  assign Black_238_io_i_pk = Black_235_io_o_p;
  assign Black_238_io_i_gk = Black_235_io_o_g;

  assign Black_240_io_i_pj = Black_438_io_o_p;
  assign Black_240_io_i_gj = Black_438_io_o_g;
  assign Black_240_io_i_pk = Black_238_io_o_p;
  assign Black_240_io_i_gk = Black_238_io_o_g;

  assign Black_242_io_i_pj = Black_463_io_o_p;
  assign Black_242_io_i_gj = Black_463_io_o_g;
  assign Black_242_io_i_pk = Black_240_io_o_p;
  assign Black_242_io_i_gk = Black_240_io_o_g;

  assign Black_246_io_i_pj = Black_486_io_o_p;
  assign Black_246_io_i_gj = Black_486_io_o_g;
  assign Black_246_io_i_pk = Black_242_io_o_p;
  assign Black_246_io_i_gk = Black_242_io_o_g;

  assign Black_248_io_i_pj = Black_514_io_o_p;
  assign Black_248_io_i_gj = Black_514_io_o_g;
  assign Black_248_io_i_pk = Black_246_io_o_p;
  assign Black_248_io_i_gk = Black_246_io_o_g;

  assign Black_251_io_i_pj = Black_524_io_o_p;
  assign Black_251_io_i_gj = Black_524_io_o_g;
  assign Black_251_io_i_pk = Black_248_io_o_p;
  assign Black_251_io_i_gk = Black_248_io_o_g;

  assign Black_253_io_i_pj = PG_275_io_o_p;
  assign Black_253_io_i_gj = PG_275_io_o_g;
  assign Black_253_io_i_pk = PG_252_io_o_p;
  assign Black_253_io_i_gk = PG_252_io_o_g;

  assign Black_254_io_i_pj = PG_297_io_o_p;
  assign Black_254_io_i_gj = PG_297_io_o_g;
  assign Black_254_io_i_pk = Black_253_io_o_p;
  assign Black_254_io_i_gk = Black_253_io_o_g;

  assign Black_257_io_i_pj = Black_320_io_o_p;
  assign Black_257_io_i_gj = Black_320_io_o_g;
  assign Black_257_io_i_pk = Black_254_io_o_p;
  assign Black_257_io_i_gk = Black_254_io_o_g;

  assign Black_258_io_i_pj = PG_375_io_o_p;
  assign Black_258_io_i_gj = PG_375_io_o_g;
  assign Black_258_io_i_pk = Black_257_io_o_p;
  assign Black_258_io_i_gk = Black_257_io_o_g;

  assign Black_263_io_i_pj = Black_396_io_o_p;
  assign Black_263_io_i_gj = Black_396_io_o_g;
  assign Black_263_io_i_pk = Black_258_io_o_p;
  assign Black_263_io_i_gk = Black_258_io_o_g;

  assign Black_274_io_i_pj = Black_472_io_o_p;
  assign Black_274_io_i_gj = Black_472_io_o_g;
  assign Black_274_io_i_pk = Black_263_io_o_p;
  assign Black_274_io_i_gk = Black_263_io_o_g;

  assign Black_276_io_i_pj = PG_297_io_o_p;
  assign Black_276_io_i_gj = PG_297_io_o_g;
  assign Black_276_io_i_pk = PG_275_io_o_p;
  assign Black_276_io_i_gk = PG_275_io_o_g;

  assign Black_280_io_i_pj = Black_321_io_o_p;
  assign Black_280_io_i_gj = Black_321_io_o_g;
  assign Black_280_io_i_pk = Black_276_io_o_p;
  assign Black_280_io_i_gk = Black_276_io_o_g;

  assign Black_289_io_i_pj = Black_400_io_o_p;
  assign Black_289_io_i_gj = Black_400_io_o_g;
  assign Black_289_io_i_pk = Black_280_io_o_p;
  assign Black_289_io_i_gk = Black_280_io_o_g;

  assign Black_296_io_i_pj = Black_506_io_o_p;
  assign Black_296_io_i_gj = Black_506_io_o_g;
  assign Black_296_io_i_pk = Black_289_io_o_p;
  assign Black_296_io_i_gk = Black_289_io_o_g;

  assign Black_298_io_i_pj = PG_318_io_o_p;
  assign Black_298_io_i_gj = PG_318_io_o_g;
  assign Black_298_io_i_pk = PG_297_io_o_p;
  assign Black_298_io_i_gk = PG_297_io_o_g;

  assign Black_317_io_i_pj = Black_356_io_o_p;
  assign Black_317_io_i_gj = Black_356_io_o_g;
  assign Black_317_io_i_pk = Black_298_io_o_p;
  assign Black_317_io_i_gk = Black_298_io_o_g;

  assign Black_319_io_i_pj = PG_338_io_o_p;
  assign Black_319_io_i_gj = PG_338_io_o_g;
  assign Black_319_io_i_pk = PG_318_io_o_p;
  assign Black_319_io_i_gk = PG_318_io_o_g;

  assign Black_320_io_i_pj = PG_357_io_o_p;
  assign Black_320_io_i_gj = PG_357_io_o_g;
  assign Black_320_io_i_pk = Black_319_io_o_p;
  assign Black_320_io_i_gk = Black_319_io_o_g;

  assign Black_321_io_i_pj = PG_375_io_o_p;
  assign Black_321_io_i_gj = PG_375_io_o_g;
  assign Black_321_io_i_pk = Black_320_io_o_p;
  assign Black_321_io_i_gk = Black_320_io_o_g;

  assign Black_337_io_i_pj = Black_407_io_o_p;
  assign Black_337_io_i_gj = Black_407_io_o_g;
  assign Black_337_io_i_pk = Black_321_io_o_p;
  assign Black_337_io_i_gk = Black_321_io_o_g;

  assign Black_340_io_i_pj = Black_358_io_o_p;
  assign Black_340_io_i_gj = Black_358_io_o_g;
  assign Black_340_io_i_pk = PG_338_io_o_p;
  assign Black_340_io_i_gk = PG_338_io_o_g;

  assign Black_352_io_i_pj = Black_403_io_o_p;
  assign Black_352_io_i_gj = Black_403_io_o_g;
  assign Black_352_io_i_pk = Black_340_io_o_p;
  assign Black_352_io_i_gk = Black_340_io_o_g;

  assign Black_356_io_i_pj = Black_521_io_o_p;
  assign Black_356_io_i_gj = Black_521_io_o_g;
  assign Black_356_io_i_pk = Black_352_io_o_p;
  assign Black_356_io_i_gk = Black_352_io_o_g;

  assign Black_358_io_i_pj = PG_375_io_o_p;
  assign Black_358_io_i_gj = PG_375_io_o_g;
  assign Black_358_io_i_pk = PG_357_io_o_p;
  assign Black_358_io_i_gk = PG_357_io_o_g;

  assign Black_363_io_i_pj = Black_396_io_o_p;
  assign Black_363_io_i_gj = Black_396_io_o_g;
  assign Black_363_io_i_pk = Black_358_io_o_p;
  assign Black_363_io_i_gk = Black_358_io_o_g;

  assign Black_374_io_i_pj = Black_472_io_o_p;
  assign Black_374_io_i_gj = Black_472_io_o_g;
  assign Black_374_io_i_pk = Black_363_io_o_p;
  assign Black_374_io_i_gk = Black_363_io_o_g;

  assign Black_391_io_i_pj = Black_407_io_o_p;
  assign Black_391_io_i_gj = Black_407_io_o_g;
  assign Black_391_io_i_pk = PG_375_io_o_p;
  assign Black_391_io_i_gk = PG_375_io_o_g;

  assign Black_393_io_i_pj = PG_408_io_o_p;
  assign Black_393_io_i_gj = PG_408_io_o_g;
  assign Black_393_io_i_pk = PG_392_io_o_p;
  assign Black_393_io_i_gk = PG_392_io_o_g;

  assign Black_394_io_i_pj = PG_423_io_o_p;
  assign Black_394_io_i_gj = PG_423_io_o_g;
  assign Black_394_io_i_pk = Black_393_io_o_p;
  assign Black_394_io_i_gk = Black_393_io_o_g;

  assign Black_395_io_i_pj = PG_437_io_o_p;
  assign Black_395_io_i_gj = PG_437_io_o_g;
  assign Black_395_io_i_pk = Black_394_io_o_p;
  assign Black_395_io_i_gk = Black_394_io_o_g;

  assign Black_396_io_i_pj = PG_450_io_o_p;
  assign Black_396_io_i_gj = PG_450_io_o_g;
  assign Black_396_io_i_pk = Black_395_io_o_p;
  assign Black_396_io_i_gk = Black_395_io_o_g;

  assign Black_398_io_i_pj = Black_463_io_o_p;
  assign Black_398_io_i_gj = Black_463_io_o_g;
  assign Black_398_io_i_pk = Black_396_io_o_p;
  assign Black_398_io_i_gk = Black_396_io_o_g;

  assign Black_399_io_i_pj = PG_483_io_o_p;
  assign Black_399_io_i_gj = PG_483_io_o_g;
  assign Black_399_io_i_pk = Black_398_io_o_p;
  assign Black_399_io_i_gk = Black_398_io_o_g;

  assign Black_400_io_i_pj = PG_492_io_o_p;
  assign Black_400_io_i_gj = PG_492_io_o_g;
  assign Black_400_io_i_pk = Black_399_io_o_p;
  assign Black_400_io_i_gk = Black_399_io_o_g;

  assign Black_403_io_i_pj = Black_502_io_o_p;
  assign Black_403_io_i_gj = Black_502_io_o_g;
  assign Black_403_io_i_pk = Black_400_io_o_p;
  assign Black_403_io_i_gk = Black_400_io_o_g;

  assign Black_407_io_i_pj = Black_521_io_o_p;
  assign Black_407_io_i_gj = Black_521_io_o_g;
  assign Black_407_io_i_pk = Black_403_io_o_p;
  assign Black_407_io_i_gk = Black_403_io_o_g;

  assign Black_414_io_i_pj = Black_428_io_o_p;
  assign Black_414_io_i_gj = Black_428_io_o_g;
  assign Black_414_io_i_pk = PG_408_io_o_p;
  assign Black_414_io_i_gk = PG_408_io_o_g;

  assign Black_416_io_i_pj = Black_493_io_o_p;
  assign Black_416_io_i_gj = Black_493_io_o_g;
  assign Black_416_io_i_pk = Black_414_io_o_p;
  assign Black_416_io_i_gk = Black_414_io_o_g;

  assign Black_422_io_i_pj = Black_512_io_o_p;
  assign Black_422_io_i_gj = Black_512_io_o_g;
  assign Black_422_io_i_pk = Black_416_io_o_p;
  assign Black_422_io_i_gk = Black_416_io_o_g;

  assign Black_428_io_i_pj = Black_441_io_o_p;
  assign Black_428_io_i_gj = Black_441_io_o_g;
  assign Black_428_io_i_pk = PG_423_io_o_p;
  assign Black_428_io_i_gk = PG_423_io_o_g;

  assign Black_432_io_i_pj = Black_495_io_o_p;
  assign Black_432_io_i_gj = Black_495_io_o_g;
  assign Black_432_io_i_pk = Black_428_io_o_p;
  assign Black_432_io_i_gk = Black_428_io_o_g;

  assign Black_436_io_i_pj = Black_521_io_o_p;
  assign Black_436_io_i_gj = Black_521_io_o_g;
  assign Black_436_io_i_pk = Black_432_io_o_p;
  assign Black_436_io_i_gk = Black_432_io_o_g;

  assign Black_438_io_i_pj = PG_450_io_o_p;
  assign Black_438_io_i_gj = PG_450_io_o_g;
  assign Black_438_io_i_pk = PG_437_io_o_p;
  assign Black_438_io_i_gk = PG_437_io_o_g;

  assign Black_441_io_i_pj = Black_464_io_o_p;
  assign Black_441_io_i_gj = Black_464_io_o_g;
  assign Black_441_io_i_pk = Black_438_io_o_p;
  assign Black_441_io_i_gk = Black_438_io_o_g;

  assign Black_448_io_i_pj = Black_498_io_o_p;
  assign Black_448_io_i_gj = Black_498_io_o_g;
  assign Black_448_io_i_pk = Black_441_io_o_p;
  assign Black_448_io_i_gk = Black_441_io_o_g;

  assign Black_449_io_i_pj = PG_527_io_o_p;
  assign Black_449_io_i_gj = PG_527_io_o_g;
  assign Black_449_io_i_pk = Black_448_io_o_p;
  assign Black_449_io_i_gk = Black_448_io_o_g;

  assign Black_451_io_i_pj = PG_462_io_o_p;
  assign Black_451_io_i_gj = PG_462_io_o_g;
  assign Black_451_io_i_pk = PG_450_io_o_p;
  assign Black_451_io_i_gk = PG_450_io_o_g;

  assign Black_458_io_i_pj = Black_479_io_o_p;
  assign Black_458_io_i_gj = Black_479_io_o_g;
  assign Black_458_io_i_pk = Black_451_io_o_p;
  assign Black_458_io_i_gk = Black_451_io_o_g;

  assign Black_461_io_i_pj = Black_524_io_o_p;
  assign Black_461_io_i_gj = Black_524_io_o_g;
  assign Black_461_io_i_pk = Black_458_io_o_p;
  assign Black_461_io_i_gk = Black_458_io_o_g;

  assign Black_463_io_i_pj = PG_473_io_o_p;
  assign Black_463_io_i_gj = PG_473_io_o_g;
  assign Black_463_io_i_pk = PG_462_io_o_p;
  assign Black_463_io_i_gk = PG_462_io_o_g;

  assign Black_464_io_i_pj = PG_483_io_o_p;
  assign Black_464_io_i_gj = PG_483_io_o_g;
  assign Black_464_io_i_pk = Black_463_io_o_p;
  assign Black_464_io_i_gk = Black_463_io_o_g;

  assign Black_467_io_i_pj = Black_494_io_o_p;
  assign Black_467_io_i_gj = Black_494_io_o_g;
  assign Black_467_io_i_pk = Black_464_io_o_p;
  assign Black_467_io_i_gk = Black_464_io_o_g;

  assign Black_469_io_i_pj = Black_514_io_o_p;
  assign Black_469_io_i_gj = Black_514_io_o_g;
  assign Black_469_io_i_pk = Black_467_io_o_p;
  assign Black_469_io_i_gk = Black_467_io_o_g;

  assign Black_472_io_i_pj = Black_524_io_o_p;
  assign Black_472_io_i_gj = Black_524_io_o_g;
  assign Black_472_io_i_pk = Black_469_io_o_p;
  assign Black_472_io_i_gk = Black_469_io_o_g;

  assign Black_478_io_i_pj = Black_487_io_o_p;
  assign Black_478_io_i_gj = Black_487_io_o_g;
  assign Black_478_io_i_pk = PG_473_io_o_p;
  assign Black_478_io_i_gk = PG_473_io_o_g;

  assign Black_479_io_i_pj = PG_518_io_o_p;
  assign Black_479_io_i_gj = PG_518_io_o_g;
  assign Black_479_io_i_pk = Black_478_io_o_p;
  assign Black_479_io_i_gk = Black_478_io_o_g;

  assign Black_482_io_i_pj = Black_524_io_o_p;
  assign Black_482_io_i_gj = Black_524_io_o_g;
  assign Black_482_io_i_pk = Black_479_io_o_p;
  assign Black_482_io_i_gk = Black_479_io_o_g;

  assign Black_486_io_i_pj = Black_494_io_o_p;
  assign Black_486_io_i_gj = Black_494_io_o_g;
  assign Black_486_io_i_pk = PG_483_io_o_p;
  assign Black_486_io_i_gk = PG_483_io_o_g;

  assign Black_487_io_i_pj = PG_513_io_o_p;
  assign Black_487_io_i_gj = PG_513_io_o_g;
  assign Black_487_io_i_pk = Black_486_io_o_p;
  assign Black_487_io_i_gk = Black_486_io_o_g;

  assign Black_491_io_i_pj = Black_521_io_o_p;
  assign Black_491_io_i_gj = Black_521_io_o_g;
  assign Black_491_io_i_pk = Black_487_io_o_p;
  assign Black_491_io_i_gk = Black_487_io_o_g;

  assign Black_493_io_i_pj = PG_500_io_o_p;
  assign Black_493_io_i_gj = PG_500_io_o_g;
  assign Black_493_io_i_pk = PG_492_io_o_p;
  assign Black_493_io_i_gk = PG_492_io_o_g;

  assign Black_494_io_i_pj = PG_507_io_o_p;
  assign Black_494_io_i_gj = PG_507_io_o_g;
  assign Black_494_io_i_pk = Black_493_io_o_p;
  assign Black_494_io_i_gk = Black_493_io_o_g;

  assign Black_495_io_i_pj = PG_513_io_o_p;
  assign Black_495_io_i_gj = PG_513_io_o_g;
  assign Black_495_io_i_pk = Black_494_io_o_p;
  assign Black_495_io_i_gk = Black_494_io_o_g;

  assign Black_497_io_i_pj = Black_519_io_o_p;
  assign Black_497_io_i_gj = Black_519_io_o_g;
  assign Black_497_io_i_pk = Black_495_io_o_p;
  assign Black_497_io_i_gk = Black_495_io_o_g;

  assign Black_498_io_i_pj = PG_525_io_o_p;
  assign Black_498_io_i_gj = PG_525_io_o_g;
  assign Black_498_io_i_pk = Black_497_io_o_p;
  assign Black_498_io_i_gk = Black_497_io_o_g;

  assign Black_499_io_i_pj = PG_527_io_o_p;
  assign Black_499_io_i_gj = PG_527_io_o_g;
  assign Black_499_io_i_pk = Black_498_io_o_p;
  assign Black_499_io_i_gk = Black_498_io_o_g;

  assign Black_502_io_i_pj = Black_508_io_o_p;
  assign Black_502_io_i_gj = Black_508_io_o_g;
  assign Black_502_io_i_pk = PG_500_io_o_p;
  assign Black_502_io_i_gk = PG_500_io_o_g;

  assign Black_503_io_i_pj = PG_518_io_o_p;
  assign Black_503_io_i_gj = PG_518_io_o_g;
  assign Black_503_io_i_pk = Black_502_io_o_p;
  assign Black_503_io_i_gk = Black_502_io_o_g;

  assign Black_506_io_i_pj = Black_524_io_o_p;
  assign Black_506_io_i_gj = Black_524_io_o_g;
  assign Black_506_io_i_pk = Black_503_io_o_p;
  assign Black_506_io_i_gk = Black_503_io_o_g;

  assign Black_508_io_i_pj = PG_513_io_o_p;
  assign Black_508_io_i_gj = PG_513_io_o_g;
  assign Black_508_io_i_pk = PG_507_io_o_p;
  assign Black_508_io_i_gk = PG_507_io_o_g;

  assign Black_512_io_i_pj = Black_521_io_o_p;
  assign Black_512_io_i_gj = Black_521_io_o_g;
  assign Black_512_io_i_pk = Black_508_io_o_p;
  assign Black_512_io_i_gk = Black_508_io_o_g;

  assign Black_514_io_i_pj = PG_518_io_o_p;
  assign Black_514_io_i_gj = PG_518_io_o_g;
  assign Black_514_io_i_pk = PG_513_io_o_p;
  assign Black_514_io_i_gk = PG_513_io_o_g;

  assign Black_515_io_i_pj = PG_522_io_o_p;
  assign Black_515_io_i_gj = PG_522_io_o_g;
  assign Black_515_io_i_pk = Black_514_io_o_p;
  assign Black_515_io_i_gk = Black_514_io_o_g;

  assign Black_517_io_i_pj = Black_526_io_o_p;
  assign Black_517_io_i_gj = Black_526_io_o_g;
  assign Black_517_io_i_pk = Black_515_io_o_p;
  assign Black_517_io_i_gk = Black_515_io_o_g;

  assign Black_519_io_i_pj = PG_522_io_o_p;
  assign Black_519_io_i_gj = PG_522_io_o_g;
  assign Black_519_io_i_pk = PG_518_io_o_p;
  assign Black_519_io_i_gk = PG_518_io_o_g;

  assign Black_521_io_i_pj = Black_526_io_o_p;
  assign Black_521_io_i_gj = Black_526_io_o_g;
  assign Black_521_io_i_pk = Black_519_io_o_p;
  assign Black_521_io_i_gk = Black_519_io_o_g;

  assign Black_523_io_i_pj = PG_525_io_o_p;
  assign Black_523_io_i_gj = PG_525_io_o_g;
  assign Black_523_io_i_pk = PG_522_io_o_p;
  assign Black_523_io_i_gk = PG_522_io_o_g;

  assign Black_524_io_i_pj = PG_527_io_o_p;
  assign Black_524_io_i_gj = PG_527_io_o_g;
  assign Black_524_io_i_pk = Black_523_io_o_p;
  assign Black_524_io_i_gk = Black_523_io_o_g;

  assign Black_526_io_i_pj = PG_527_io_o_p;
  assign Black_526_io_i_gj = PG_527_io_o_g;
  assign Black_526_io_i_pk = PG_525_io_o_p;
  assign Black_526_io_i_gk = PG_525_io_o_g;

endmodule
module MultTop (
    input clock,
  input reset,

  input [15:0] multiplicand,
  input [15:0] multiplier,
  output [31:0] product
);
  wire [0:0] pp_0;
  wire [1:0] pp_1;
  wire [2:0] pp_2;
  wire [3:0] pp_3;
  wire [4:0] pp_4;
  wire [5:0] pp_5;
  wire [6:0] pp_6;
  wire [7:0] pp_7;
  wire [8:0] pp_8;
  wire [9:0] pp_9;
  wire [10:0] pp_10;
  wire [11:0] pp_11;
  wire [12:0] pp_12;
  wire [13:0] pp_13;
  wire [14:0] pp_14;
  wire [15:0] pp_15;
  wire [14:0] pp_16;
  wire [13:0] pp_17;
  wire [12:0] pp_18;
  wire [11:0] pp_19;
  wire [10:0] pp_20;
  wire [9:0] pp_21;
  wire [8:0] pp_22;
  wire [7:0] pp_23;
  wire [6:0] pp_24;
  wire [5:0] pp_25;
  wire [4:0] pp_26;
  wire [3:0] pp_27;
  wire [2:0] pp_28;
  wire [1:0] pp_29;
  wire [0:0] pp_30;
  wire [31:0] augend;
  wire [31:0] addend;

  PartialProductGenerator pp_gen(
    .pp_0(pp_0),
    .pp_1(pp_1),
    .pp_2(pp_2),
    .pp_3(pp_3),
    .pp_4(pp_4),
    .pp_5(pp_5),
    .pp_6(pp_6),
    .pp_7(pp_7),
    .pp_8(pp_8),
    .pp_9(pp_9),
    .pp_10(pp_10),
    .pp_11(pp_11),
    .pp_12(pp_12),
    .pp_13(pp_13),
    .pp_14(pp_14),
    .pp_15(pp_15),
    .pp_16(pp_16),
    .pp_17(pp_17),
    .pp_18(pp_18),
    .pp_19(pp_19),
    .pp_20(pp_20),
    .pp_21(pp_21),
    .pp_22(pp_22),
    .pp_23(pp_23),
    .pp_24(pp_24),
    .pp_25(pp_25),
    .pp_26(pp_26),
    .pp_27(pp_27),
    .pp_28(pp_28),
    .pp_29(pp_29),
    .pp_30(pp_30),
    .multiplicand(multiplicand),
    .multiplier(multiplier)
  );

  CompressorTree comp_tree(
    .io_pp_0(pp_0),
    .io_pp_1(pp_1),
    .io_pp_2(pp_2),
    .io_pp_3(pp_3),
    .io_pp_4(pp_4),
    .io_pp_5(pp_5),
    .io_pp_6(pp_6),
    .io_pp_7(pp_7),
    .io_pp_8(pp_8),
    .io_pp_9(pp_9),
    .io_pp_10(pp_10),
    .io_pp_11(pp_11),
    .io_pp_12(pp_12),
    .io_pp_13(pp_13),
    .io_pp_14(pp_14),
    .io_pp_15(pp_15),
    .io_pp_16(pp_16),
    .io_pp_17(pp_17),
    .io_pp_18(pp_18),
    .io_pp_19(pp_19),
    .io_pp_20(pp_20),
    .io_pp_21(pp_21),
    .io_pp_22(pp_22),
    .io_pp_23(pp_23),
    .io_pp_24(pp_24),
    .io_pp_25(pp_25),
    .io_pp_26(pp_26),
    .io_pp_27(pp_27),
    .io_pp_28(pp_28),
    .io_pp_29(pp_29),
    .io_pp_30(pp_30),
    .io_augend(augend),
    .io_addend(addend)
  );

  CarryPropagateAdder final_adder(
    .io_augend(augend),
    .io_addend(addend),
    .io_outs(product)
  );

endmodule
