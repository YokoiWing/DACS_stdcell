# BSD 3-Clause License
# 
# Copyright 2020 Lawrence T. Clark, Vinay Vashishtha, or Arizona State
# University
# 
# Redistribution and use in source and binary forms, with or without
# modification, are permitted provided that the following conditions are met:
# 
# 1. Redistributions of source code must retain the above copyright notice,
# this list of conditions and the following disclaimer.
# 
# 2. Redistributions in binary form must reproduce the above copyright
# notice, this list of conditions and the following disclaimer in the
# documentation and/or other materials provided with the distribution.
# 
# 3. Neither the name of the copyright holder nor the names of its
# contributors may be used to endorse or promote products derived from this
# software without specific prior written permission.
# 
# THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
# AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
# IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
# ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
# LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
# CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
# SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
# INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
# CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
# ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
# POSSIBILITY OF SUCH DAMAGE.

VERSION 5.8 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 


SITE asap7sc7p5t 
 CLASS CORE ; 
 SIZE 0.216 BY 1.08 ; 
 SYMMETRY Y ; 
END asap7sc7p5t 


MACRO A2O1A1Ixp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN A2O1A1Ixp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.324 1.008 0.76 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.856 0.86 1.224 0.932 ; 
        RECT 1.152 0.148 1.224 0.932 ; 
        RECT 1.048 0.148 1.224 0.22 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 0.92 0.18 ; 
      RECT 0.16 0.9 0.704 0.972 ; 
  END 
END A2O1A1Ixp33_ASAP7_75t_R 


MACRO A2O1A1O1Ixp25_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN A2O1A1O1Ixp25_ASAP7_75t_R 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.508 1.656 0.58 ; 
        RECT 1.368 0.28 1.44 0.8 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.944 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.692 0.9 1.872 0.972 ; 
        RECT 1.8 0.108 1.872 0.972 ; 
        RECT 1.044 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.828 0.9 1.548 0.972 ; 
      RECT 0.16 0.108 0.9 0.18 ; 
      RECT 0.16 0.9 0.684 0.972 ; 
  END 
END A2O1A1O1Ixp25_ASAP7_75t_R 


MACRO AND2x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x2_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.336 0.576 ; 
        RECT 0.072 0.136 0.144 0.944 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.9 1.224 0.972 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
        RECT 0.828 0.108 1.224 0.18 ; 
        RECT 0.828 0.736 0.9 0.972 ; 
        RECT 0.828 0.108 0.9 0.344 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.9 0.72 0.972 ; 
      RECT 0.648 0.108 0.72 0.972 ; 
      RECT 0.648 0.504 0.812 0.576 ; 
      RECT 0.28 0.108 0.352 0.344 ; 
      RECT 0.28 0.108 0.72 0.18 ; 
  END 
END AND2x2_ASAP7_75t_R 


MACRO AND2x4_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x4_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.112 1.008 0.6 ; 
        RECT 0.288 0.112 1.008 0.184 ; 
        RECT 0.288 0.112 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.428 0.576 0.8 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.9 1.872 0.972 ; 
        RECT 1.8 0.108 1.872 0.972 ; 
        RECT 1.24 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.9 0.924 0.972 ; 
      RECT 0.72 0.256 0.792 0.972 ; 
      RECT 0.716 0.728 1.224 0.8 ; 
      RECT 1.152 0.484 1.224 0.8 ; 
      RECT 0.46 0.256 0.792 0.328 ; 
  END 
END AND2x4_ASAP7_75t_R 


MACRO AND2x6_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND2x6_ASAP7_75t_R 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.112 1.008 0.6 ; 
        RECT 0.288 0.112 1.008 0.184 ; 
        RECT 0.288 0.112 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.428 0.576 0.8 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.592 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.9 2.216 0.972 ; 
        RECT 1.24 0.108 2.216 0.18 ; 
        RECT 1.8 0.108 1.872 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.9 0.924 0.972 ; 
      RECT 0.72 0.256 0.792 0.972 ; 
      RECT 0.716 0.728 1.224 0.8 ; 
      RECT 1.152 0.484 1.224 0.8 ; 
      RECT 0.46 0.256 0.792 0.328 ; 
  END 
END AND2x6_ASAP7_75t_R 


MACRO AND3x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND3x1_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.732 1.224 0.804 ; 
        RECT 1.152 0.304 1.224 0.804 ; 
        RECT 1.044 0.304 1.224 0.376 ; 
        RECT 1.044 0.732 1.116 0.94 ; 
        RECT 1.044 0.136 1.116 0.376 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.936 0.972 ; 
      RECT 0.864 0.108 0.936 0.972 ; 
      RECT 0.864 0.504 1.052 0.576 ; 
      RECT 0.16 0.108 0.936 0.18 ; 
  END 
END AND3x1_ASAP7_75t_R 


MACRO AND3x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND3x2_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.9 1.44 0.972 ; 
        RECT 1.368 0.108 1.44 0.972 ; 
        RECT 1.044 0.108 1.44 0.18 ; 
        RECT 1.044 0.736 1.116 0.972 ; 
        RECT 1.044 0.108 1.116 0.344 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.936 0.972 ; 
      RECT 0.864 0.108 0.936 0.972 ; 
      RECT 0.864 0.504 1.136 0.576 ; 
      RECT 0.16 0.108 0.936 0.18 ; 
  END 
END AND3x2_ASAP7_75t_R 


MACRO AND3x4_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND3x4_ASAP7_75t_R 0 0 ; 
  SIZE 3.024 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.448 0.756 2.596 0.828 ; 
        RECT 2.448 0.396 2.596 0.468 ; 
        RECT 2.448 0.396 2.52 0.828 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.756 2.164 0.828 ; 
        RECT 2.016 0.396 2.164 0.468 ; 
        RECT 2.016 0.396 2.088 0.828 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.8 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.024 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.92 0.972 ; 
        RECT 0.072 0.108 0.92 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.04 0.9 2.984 0.972 ; 
      RECT 2.912 0.108 2.984 0.972 ; 
      RECT 1.04 0.168 1.112 0.972 ; 
      RECT 0.872 0.504 1.112 0.576 ; 
      RECT 2.536 0.108 2.984 0.18 ; 
      RECT 1.888 0.252 2.804 0.324 ; 
      RECT 1.24 0.108 2.216 0.18 ; 
  END 
END AND3x4_ASAP7_75t_R 


MACRO AND4x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND4x1_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.136 0.576 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.136 0.792 0.8 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.136 1.008 0.656 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.196 0.9 1.44 0.972 ; 
        RECT 1.368 0.108 1.44 0.972 ; 
        RECT 1.24 0.108 1.44 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.072 0.9 1.008 0.972 ; 
      RECT 0.936 0.756 1.008 0.972 ; 
      RECT 0.072 0.108 0.144 0.972 ; 
      RECT 0.936 0.756 1.224 0.828 ; 
      RECT 1.152 0.48 1.224 0.828 ; 
      RECT 0.072 0.108 0.34 0.18 ; 
  END 
END AND4x1_ASAP7_75t_R 


MACRO AND4x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND4x2_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.136 1.224 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.136 1.008 0.8 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.136 0.792 0.656 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.488 0.972 ; 
        RECT 0.072 0.108 0.488 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.612 0.9 1.656 0.972 ; 
      RECT 1.584 0.108 1.656 0.972 ; 
      RECT 0.612 0.756 0.684 0.972 ; 
      RECT 0.396 0.756 0.684 0.828 ; 
      RECT 0.396 0.476 0.468 0.828 ; 
      RECT 1.456 0.108 1.656 0.18 ; 
  END 
END AND4x2_ASAP7_75t_R 


MACRO AND5x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND5x1_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.136 0.576 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.136 0.792 0.8 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.136 1.008 0.8 ; 
    END 
  END D 
  PIN E 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.136 1.224 0.656 ; 
    END 
  END E 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.396 0.9 1.656 0.972 ; 
        RECT 1.584 0.108 1.656 0.972 ; 
        RECT 1.4 0.108 1.656 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.072 0.9 1.224 0.972 ; 
      RECT 1.152 0.756 1.224 0.972 ; 
      RECT 0.072 0.108 0.144 0.972 ; 
      RECT 1.152 0.756 1.44 0.828 ; 
      RECT 1.368 0.464 1.44 0.828 ; 
      RECT 0.072 0.108 0.28 0.18 ; 
  END 
END AND5x1_ASAP7_75t_R 


MACRO AND5x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AND5x2_ASAP7_75t_R 0 0 ; 
  SIZE 4.32 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.88 0.756 3.028 0.828 ; 
        RECT 2.88 0.396 3.028 0.468 ; 
        RECT 2.88 0.396 2.952 0.828 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.372 0.756 2.52 0.828 ; 
        RECT 2.448 0.396 2.52 0.828 ; 
        RECT 2.372 0.396 2.52 0.468 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.756 1.948 0.828 ; 
        RECT 1.8 0.396 1.948 0.468 ; 
        RECT 1.8 0.396 1.872 0.828 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.076 0.756 1.224 0.828 ; 
        RECT 1.152 0.396 1.224 0.828 ; 
        RECT 1.076 0.396 1.224 0.468 ; 
    END 
  END D 
  PIN E 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.136 0.144 0.944 ; 
    END 
  END E 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.32 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.32 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.832 0.9 4.248 0.972 ; 
        RECT 4.176 0.108 4.248 0.972 ; 
        RECT 3.832 0.108 4.248 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.592 0.9 3.6 0.972 ; 
      RECT 3.528 0.108 3.6 0.972 ; 
      RECT 3.528 0.504 3.768 0.576 ; 
      RECT 2.968 0.108 3.6 0.18 ; 
      RECT 2.32 0.252 3.296 0.324 ; 
      RECT 1.672 0.108 2.648 0.18 ; 
      RECT 1.024 0.252 2 0.324 ; 
      RECT 0.376 0.108 1.352 0.18 ; 
  END 
END AND5x2_ASAP7_75t_R 


MACRO AO211x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO211x2_ASAP7_75t_R 0 0 ; 
  SIZE 3.456 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.828 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.504 0.812 0.576 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.504 1.244 0.576 ; 
        RECT 0.86 0.756 1.008 0.828 ; 
        RECT 0.936 0.252 1.008 0.828 ; 
        RECT 0.86 0.252 1.008 0.324 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.612 2.164 0.684 ; 
        RECT 2.016 0.252 2.088 0.684 ; 
        RECT 1.94 0.252 2.088 0.324 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.456 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.456 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.968 0.9 3.384 0.972 ; 
        RECT 3.312 0.108 3.384 0.972 ; 
        RECT 2.968 0.108 3.384 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.104 0.9 2.736 0.972 ; 
      RECT 2.664 0.108 2.736 0.972 ; 
      RECT 2.664 0.5 2.972 0.572 ; 
      RECT 0.376 0.108 2.736 0.18 ; 
      RECT 1.24 0.756 2.432 0.828 ; 
      RECT 0.16 0.9 1.572 0.972 ; 
  END 
END AO211x2_ASAP7_75t_R 


MACRO AO21x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21x1_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.136 0.144 0.828 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.656 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.92 0.9 1.18 0.972 ; 
        RECT 1.108 0.152 1.18 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.756 1.008 0.828 ; 
      RECT 0.936 0.108 1.008 0.828 ; 
      RECT 0.592 0.108 1.008 0.18 ; 
      RECT 0.16 0.9 0.704 0.972 ; 
  END 
END AO21x1_ASAP7_75t_R 


MACRO AO21x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO21x2_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.136 0.144 0.828 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.656 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.92 0.9 1.332 0.972 ; 
        RECT 1.26 0.276 1.332 0.972 ; 
        RECT 1.104 0.276 1.332 0.348 ; 
        RECT 1.104 0.152 1.176 0.348 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.756 1.008 0.828 ; 
      RECT 0.936 0.108 1.008 0.828 ; 
      RECT 0.592 0.108 1.008 0.18 ; 
      RECT 0.16 0.9 0.704 0.972 ; 
  END 
END AO21x2_ASAP7_75t_R 


MACRO AO221x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO221x1_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.656 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.656 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.888 0.9 2.088 0.972 ; 
        RECT 2.016 0.108 2.088 0.972 ; 
        RECT 1.836 0.108 2.088 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.072 0.756 0.504 0.828 ; 
      RECT 0.072 0.108 0.144 0.828 ; 
      RECT 1.584 0.504 1.896 0.576 ; 
      RECT 1.584 0.108 1.656 0.576 ; 
      RECT 0.072 0.108 1.656 0.18 ; 
      RECT 0.8 0.756 1.356 0.828 ; 
      RECT 0.156 0.9 0.704 0.972 ; 
  END 
END AO221x1_ASAP7_75t_R 


MACRO AO221x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO221x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.656 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.656 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.888 0.9 2.196 0.972 ; 
        RECT 2.124 0.108 2.196 0.972 ; 
        RECT 1.836 0.108 2.196 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.072 0.756 0.504 0.828 ; 
      RECT 0.072 0.108 0.144 0.828 ; 
      RECT 1.584 0.504 1.896 0.576 ; 
      RECT 1.584 0.108 1.656 0.576 ; 
      RECT 0.072 0.108 1.656 0.18 ; 
      RECT 0.8 0.756 1.356 0.828 ; 
      RECT 0.156 0.9 0.704 0.972 ; 
  END 
END AO221x2_ASAP7_75t_R 


MACRO AO222x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO222x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.28 1.872 0.8 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.656 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.656 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.592 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.104 0.9 2.52 0.972 ; 
        RECT 2.448 0.108 2.52 0.972 ; 
        RECT 2.124 0.108 2.52 0.18 ; 
        RECT 2.124 0.108 2.196 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.036 0.756 0.488 0.828 ; 
      RECT 0.036 0.108 0.108 0.828 ; 
      RECT 1.944 0.504 2.216 0.576 ; 
      RECT 1.944 0.108 2.016 0.576 ; 
      RECT 0.036 0.108 2.016 0.18 ; 
      RECT 1.368 0.9 1.872 0.972 ; 
      RECT 1.368 0.756 1.44 0.972 ; 
      RECT 0.808 0.756 1.44 0.828 ; 
      RECT 0.16 0.9 1.136 0.972 ; 
  END 
END AO222x2_ASAP7_75t_R 


MACRO AO22x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO22x1_ASAP7_75t_R 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.828 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.252 1.148 0.324 ; 
        RECT 0.936 0.252 1.008 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.944 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.9 1.872 0.972 ; 
        RECT 1.8 0.108 1.872 0.972 ; 
        RECT 1.672 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.808 0.756 1.44 0.828 ; 
      RECT 1.368 0.108 1.44 0.828 ; 
      RECT 1.368 0.504 1.676 0.576 ; 
      RECT 0.428 0.108 1.44 0.18 ; 
      RECT 0.16 0.9 1.136 0.972 ; 
  END 
END AO22x1_ASAP7_75t_R 


MACRO AO22x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO22x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.828 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.252 1.148 0.324 ; 
        RECT 0.936 0.252 1.008 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.9 2.088 0.972 ; 
        RECT 2.016 0.108 2.088 0.972 ; 
        RECT 1.672 0.108 2.088 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.808 0.756 1.44 0.828 ; 
      RECT 1.368 0.108 1.44 0.828 ; 
      RECT 1.368 0.504 1.676 0.576 ; 
      RECT 0.428 0.108 1.44 0.18 ; 
      RECT 0.16 0.9 1.136 0.972 ; 
  END 
END AO22x2_ASAP7_75t_R 


MACRO AO31x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO31x2_ASAP7_75t_R 0 0 ; 
  SIZE 3.456 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.232 0.396 2.304 0.596 ; 
        RECT 2.016 0.396 2.304 0.468 ; 
        RECT 1.94 0.612 2.088 0.684 ; 
        RECT 2.016 0.396 2.088 0.684 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.396 1.656 0.596 ; 
        RECT 1.152 0.396 1.656 0.468 ; 
        RECT 1.152 0.612 1.3 0.684 ; 
        RECT 1.152 0.28 1.224 0.684 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.756 0.236 0.828 ; 
        RECT 0.072 0.108 0.236 0.18 ; 
        RECT 0.072 0.108 0.144 0.828 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.504 0.812 0.576 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.456 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.456 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.964 0.9 3.384 0.972 ; 
        RECT 3.312 0.108 3.384 0.972 ; 
        RECT 2.968 0.108 3.384 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.448 0.9 2.736 0.972 ; 
      RECT 2.664 0.108 2.736 0.972 ; 
      RECT 2.448 0.756 2.52 0.972 ; 
      RECT 0.796 0.756 2.52 0.828 ; 
      RECT 0.936 0.252 1.008 0.828 ; 
      RECT 2.664 0.504 3.188 0.576 ; 
      RECT 0.8 0.252 1.008 0.324 ; 
      RECT 2.104 0.108 2.736 0.18 ; 
      RECT 1.456 0.252 2.432 0.324 ; 
      RECT 0.16 0.9 2.216 0.972 ; 
      RECT 0.376 0.108 1.788 0.18 ; 
  END 
END AO31x2_ASAP7_75t_R 


MACRO AO322x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO322x2_ASAP7_75t_R 0 0 ; 
  SIZE 3.24 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.972 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.612 1.3 0.684 ; 
        RECT 1.152 0.252 1.3 0.324 ; 
        RECT 1.152 0.252 1.224 0.684 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.28 1.872 0.656 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.252 2.164 0.324 ; 
        RECT 2.016 0.252 2.088 0.656 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.24 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.24 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.536 0.9 3.168 0.972 ; 
        RECT 3.096 0.108 3.168 0.972 ; 
        RECT 2.536 0.108 3.168 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.584 0.756 2.304 0.828 ; 
      RECT 2.232 0.504 2.304 0.828 ; 
      RECT 1.584 0.108 1.656 0.828 ; 
      RECT 2.232 0.504 2.972 0.576 ; 
      RECT 0.16 0.108 1.784 0.18 ; 
      RECT 0.376 0.9 0.792 0.972 ; 
      RECT 0.72 0.756 0.792 0.972 ; 
      RECT 0.72 0.756 1.352 0.828 ; 
      RECT 1.024 0.9 2 0.972 ; 
  END 
END AO322x2_ASAP7_75t_R 


MACRO AO32x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO32x1_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.272 0.972 ; 
        RECT 0.072 0.252 0.252 0.324 ; 
        RECT 0.18 0.136 0.252 0.324 ; 
        RECT 0.072 0.252 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.24 0.756 1.656 0.828 ; 
      RECT 1.584 0.108 1.656 0.828 ; 
      RECT 0.248 0.504 0.432 0.576 ; 
      RECT 0.36 0.108 0.432 0.576 ; 
      RECT 0.36 0.108 1.656 0.18 ; 
      RECT 0.592 0.9 1.568 0.972 ; 
  END 
END AO32x1_ASAP7_75t_R 


MACRO AO32x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO32x2_ASAP7_75t_R 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.756 1.32 0.828 ; 
        RECT 1.152 0.28 1.224 0.828 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.656 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.944 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.488 0.972 ; 
        RECT 0.072 0.272 0.468 0.344 ; 
        RECT 0.396 0.148 0.468 0.344 ; 
        RECT 0.072 0.272 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.456 0.756 1.872 0.828 ; 
      RECT 1.8 0.108 1.872 0.828 ; 
      RECT 0.372 0.504 0.648 0.576 ; 
      RECT 0.576 0.108 0.648 0.576 ; 
      RECT 0.576 0.108 1.872 0.18 ; 
      RECT 0.808 0.9 1.784 0.972 ; 
  END 
END AO32x2_ASAP7_75t_R 


MACRO AO331x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO331x1_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.656 ; 
    END 
  END B3 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.28 1.872 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.324 0.18 ; 
        RECT 0.072 0.9 0.272 0.972 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.884 0.9 2.088 0.972 ; 
      RECT 2.016 0.108 2.088 0.972 ; 
      RECT 0.288 0.252 0.36 0.608 ; 
      RECT 0.288 0.252 0.576 0.324 ; 
      RECT 0.504 0.108 0.576 0.324 ; 
      RECT 0.504 0.108 2.088 0.18 ; 
      RECT 1.232 0.756 1.788 0.828 ; 
      RECT 0.584 0.9 1.572 0.972 ; 
  END 
END AO331x1_ASAP7_75t_R 


MACRO AO331x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO331x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.656 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.28 1.872 0.656 ; 
    END 
  END B3 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.28 2.088 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.108 0.54 0.18 ; 
        RECT 0.288 0.9 0.488 0.972 ; 
        RECT 0.288 0.108 0.36 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.1 0.9 2.304 0.972 ; 
      RECT 2.232 0.108 2.304 0.972 ; 
      RECT 0.504 0.252 0.576 0.608 ; 
      RECT 0.504 0.252 0.792 0.324 ; 
      RECT 0.72 0.108 0.792 0.324 ; 
      RECT 0.72 0.108 2.304 0.18 ; 
      RECT 1.448 0.756 2.004 0.828 ; 
      RECT 0.8 0.9 1.788 0.972 ; 
  END 
END AO331x2_ASAP7_75t_R 


MACRO AO332x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO332x1_ASAP7_75t_R 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.656 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.28 2.088 0.656 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.28 1.872 0.656 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.376 0.18 ; 
        RECT 0.072 0.9 0.272 0.972 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.884 0.756 2.304 0.828 ; 
      RECT 2.232 0.108 2.304 0.828 ; 
      RECT 0.288 0.252 0.36 0.604 ; 
      RECT 0.288 0.252 0.576 0.324 ; 
      RECT 0.504 0.108 0.576 0.324 ; 
      RECT 0.504 0.108 2.304 0.18 ; 
      RECT 0.584 0.9 1.008 0.972 ; 
      RECT 0.936 0.756 1.008 0.972 ; 
      RECT 0.936 0.756 1.572 0.828 ; 
      RECT 1.232 0.9 2.224 0.972 ; 
  END 
END AO332x1_ASAP7_75t_R 


MACRO AO332x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO332x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.656 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.656 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.28 1.872 0.656 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.232 0.28 2.304 0.656 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.28 2.088 0.656 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.592 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.592 0.18 ; 
        RECT 0.072 0.9 0.488 0.972 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.1 0.756 2.52 0.828 ; 
      RECT 2.448 0.108 2.52 0.828 ; 
      RECT 0.504 0.252 0.576 0.604 ; 
      RECT 0.504 0.252 0.792 0.324 ; 
      RECT 0.72 0.108 0.792 0.324 ; 
      RECT 0.72 0.108 2.52 0.18 ; 
      RECT 0.8 0.9 1.224 0.972 ; 
      RECT 1.152 0.756 1.224 0.972 ; 
      RECT 1.152 0.756 1.788 0.828 ; 
      RECT 1.448 0.9 2.44 0.972 ; 
  END 
END AO332x2_ASAP7_75t_R 


MACRO AO333x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO333x1_ASAP7_75t_R 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.656 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.232 0.28 2.304 0.656 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.28 2.088 0.656 ; 
    END 
  END C2 
  PIN C3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.28 1.872 0.656 ; 
    END 
  END C3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.592 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.324 0.18 ; 
        RECT 0.072 0.9 0.276 0.972 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.884 0.9 2.52 0.972 ; 
      RECT 2.448 0.108 2.52 0.972 ; 
      RECT 0.288 0.252 0.36 0.608 ; 
      RECT 0.288 0.252 0.576 0.324 ; 
      RECT 0.504 0.108 0.576 0.324 ; 
      RECT 0.504 0.108 2.52 0.18 ; 
      RECT 1.24 0.756 2.304 0.828 ; 
      RECT 0.592 0.9 1.58 0.972 ; 
  END 
END AO333x1_ASAP7_75t_R 


MACRO AO333x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO333x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.808 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.28 1.872 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.656 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.448 0.28 2.52 0.656 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.232 0.28 2.304 0.656 ; 
    END 
  END C2 
  PIN C3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.28 2.088 0.656 ; 
    END 
  END C3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.808 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.808 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.488 0.972 ; 
        RECT 0.072 0.324 0.468 0.396 ; 
        RECT 0.396 0.18 0.468 0.396 ; 
        RECT 0.072 0.324 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.1 0.9 2.736 0.972 ; 
      RECT 2.664 0.108 2.736 0.972 ; 
      RECT 0.268 0.504 0.648 0.576 ; 
      RECT 0.576 0.108 0.648 0.576 ; 
      RECT 0.576 0.108 2.736 0.18 ; 
      RECT 1.456 0.756 2.52 0.828 ; 
      RECT 0.808 0.9 1.796 0.972 ; 
  END 
END AO333x2_ASAP7_75t_R 


MACRO AO33x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AO33x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.656 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.28 1.872 0.656 ; 
    END 
  END B3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.488 0.972 ; 
        RECT 0.072 0.272 0.468 0.344 ; 
        RECT 0.396 0.148 0.468 0.344 ; 
        RECT 0.072 0.272 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.444 0.756 2.088 0.828 ; 
      RECT 2.016 0.108 2.088 0.828 ; 
      RECT 0.268 0.504 0.648 0.576 ; 
      RECT 0.576 0.108 0.648 0.576 ; 
      RECT 0.576 0.108 2.088 0.18 ; 
      RECT 0.796 0.9 1.796 0.972 ; 
  END 
END AO33x2_ASAP7_75t_R 


MACRO AOI211x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI211x1_ASAP7_75t_R 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.504 0.916 0.576 ; 
        RECT 0.72 0.756 0.892 0.828 ; 
        RECT 0.72 0.252 0.88 0.324 ; 
        RECT 0.72 0.252 0.792 0.828 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.492 0.576 ; 
        RECT 0.072 0.136 0.144 0.944 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.612 1.768 0.684 ; 
        RECT 1.584 0.252 1.768 0.324 ; 
        RECT 1.584 0.252 1.656 0.684 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.504 2.216 0.576 ; 
        RECT 2.016 0.252 2.2 0.324 ; 
        RECT 2.016 0.252 2.088 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.592 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.076 0.756 2.52 0.828 ; 
        RECT 2.448 0.108 2.52 0.828 ; 
        RECT 0.364 0.108 2.52 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.364 0.9 1.224 0.972 ; 
      RECT 1.152 0.756 1.224 0.972 ; 
      RECT 1.152 0.756 1.796 0.828 ; 
      RECT 1.444 0.9 2.432 0.972 ; 
  END 
END AOI211x1_ASAP7_75t_R 


MACRO AOI211xp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI211xp5_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.656 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.36 0.576 ; 
        RECT 0.072 0.28 0.144 0.8 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.756 1.224 0.828 ; 
        RECT 1.152 0.108 1.224 0.828 ; 
        RECT 0.16 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.704 0.972 ; 
  END 
END AOI211xp5_ASAP7_75t_R 


MACRO AOI21x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21x1_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.252 1.224 0.656 ; 
        RECT 0.504 0.252 1.224 0.324 ; 
        RECT 0.504 0.252 0.576 0.656 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.76 0.5 1.024 0.572 ; 
        RECT 0.76 0.396 0.908 0.684 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.756 1.44 0.828 ; 
        RECT 1.368 0.464 1.44 0.828 ; 
        RECT 0.288 0.28 0.36 0.828 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.476 0.9 1.656 0.972 ; 
        RECT 1.584 0.108 1.656 0.972 ; 
        RECT 0.072 0.108 1.656 0.18 ; 
        RECT 0.072 0.9 0.252 0.972 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.9 1.332 0.972 ; 
  END 
END AOI21x1_ASAP7_75t_R 


MACRO AOI21xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.08 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.5 0.38 0.572 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.828 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.08 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.9 1.008 0.972 ; 
        RECT 0.936 0.108 1.008 0.972 ; 
        RECT 0.428 0.108 1.008 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.684 0.972 ; 
  END 
END AOI21xp33_ASAP7_75t_R 


MACRO AOI21xp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI21xp5_ASAP7_75t_R 0 0 ; 
  SIZE 1.08 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.5 0.38 0.572 ; 
        RECT 0.072 0.136 0.144 0.8 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.08 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.9 1.008 0.972 ; 
        RECT 0.936 0.108 1.008 0.972 ; 
        RECT 0.568 0.108 1.008 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.684 0.972 ; 
  END 
END AOI21xp5_ASAP7_75t_R 


MACRO AOI221x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI221x1_ASAP7_75t_R 0 0 ; 
  SIZE 3.024 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.612 0.868 0.684 ; 
        RECT 0.72 0.108 0.792 0.684 ; 
        RECT 0.644 0.108 0.792 0.18 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.504 0.596 0.576 ; 
        RECT 0.212 0.612 0.36 0.684 ; 
        RECT 0.288 0.108 0.36 0.684 ; 
        RECT 0.212 0.108 0.36 0.18 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.324 1.3 0.396 ; 
        RECT 1.076 0.612 1.224 0.684 ; 
        RECT 1.152 0.324 1.224 0.684 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.612 1.948 0.684 ; 
        RECT 1.8 0.324 1.872 0.684 ; 
        RECT 1.564 0.504 1.872 0.576 ; 
        RECT 1.724 0.324 1.872 0.396 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.232 0.504 2.544 0.576 ; 
        RECT 2.156 0.756 2.304 0.828 ; 
        RECT 2.232 0.324 2.304 0.828 ; 
        RECT 2.156 0.324 2.304 0.396 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.024 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.536 0.756 2.952 0.828 ; 
        RECT 2.88 0.18 2.952 0.828 ; 
        RECT 1.024 0.18 2.952 0.252 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.24 0.9 2.864 0.972 ; 
      RECT 0.16 0.756 2 0.828 ; 
  END 
END AOI221x1_ASAP7_75t_R 


MACRO AOI221xp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI221xp5_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.136 1.224 0.656 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.656 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.92 0.18 ; 
        RECT 0.072 0.756 0.492 0.828 ; 
        RECT 0.072 0.108 0.144 0.828 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.804 0.756 1.356 0.828 ; 
      RECT 0.16 0.9 0.704 0.972 ; 
  END 
END AOI221xp5_ASAP7_75t_R 


MACRO AOI222xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI222xp33_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.656 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.656 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.8 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.136 1.872 0.8 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 1.596 0.18 ; 
        RECT 0.072 0.756 0.488 0.828 ; 
        RECT 0.072 0.108 0.144 0.828 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.368 0.9 1.872 0.972 ; 
      RECT 1.368 0.756 1.44 0.972 ; 
      RECT 0.808 0.756 1.44 0.828 ; 
      RECT 0.16 0.9 1.136 0.972 ; 
  END 
END AOI222xp33_ASAP7_75t_R 


MACRO AOI22x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI22x1_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.612 1.516 0.684 ; 
        RECT 1.368 0.396 1.516 0.468 ; 
        RECT 1.368 0.396 1.44 0.684 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.724 0.612 1.872 0.684 ; 
        RECT 1.8 0.252 1.872 0.684 ; 
        RECT 1.152 0.252 1.872 0.324 ; 
        RECT 1.152 0.252 1.224 0.608 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.644 0.756 0.792 0.828 ; 
        RECT 0.72 0.396 0.792 0.828 ; 
        RECT 0.644 0.396 0.792 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.252 1.008 0.616 ; 
        RECT 0.288 0.252 1.008 0.324 ; 
        RECT 0.288 0.756 0.436 0.828 ; 
        RECT 0.288 0.252 0.36 0.828 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.236 0.756 2.088 0.828 ; 
        RECT 2.016 0.108 2.088 0.828 ; 
        RECT 0.152 0.108 2.088 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 2 0.972 ; 
  END 
END AOI22x1_ASAP7_75t_R 


MACRO AOI22xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI22xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.136 0.36 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.756 1.224 0.828 ; 
        RECT 1.152 0.108 1.224 0.828 ; 
        RECT 0.592 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 1.136 0.972 ; 
  END 
END AOI22xp33_ASAP7_75t_R 


MACRO AOI22xp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI22xp5_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.828 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.28 0.576 0.828 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.756 1.224 0.828 ; 
        RECT 1.152 0.108 1.224 0.828 ; 
        RECT 0.592 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 1.136 0.972 ; 
  END 
END AOI22xp5_ASAP7_75t_R 


MACRO AOI311xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI311xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.136 0.576 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.136 0.144 0.944 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.8 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.9 1.44 0.972 ; 
        RECT 1.368 0.108 1.44 0.972 ; 
        RECT 0.792 0.108 1.44 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.9 0.936 0.972 ; 
  END 
END AOI311xp33_ASAP7_75t_R 


MACRO AOI31xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI31xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.136 0.576 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.136 0.36 0.8 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.756 1.224 0.828 ; 
        RECT 1.152 0.108 1.224 0.828 ; 
        RECT 0.804 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.372 0.9 0.92 0.972 ; 
  END 
END AOI31xp33_ASAP7_75t_R 


MACRO AOI31xp67_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI31xp67_ASAP7_75t_R 0 0 ; 
  SIZE 2.808 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.664 0.28 2.736 0.8 ; 
        RECT 2.212 0.504 2.736 0.576 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.504 1.676 0.576 ; 
        RECT 1.152 0.252 1.3 0.324 ; 
        RECT 1.152 0.252 1.224 0.656 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.756 0.236 0.828 ; 
        RECT 0.072 0.108 0.236 0.18 ; 
        RECT 0.072 0.108 0.144 0.828 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.504 0.812 0.576 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.808 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.808 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.34 0.9 2.652 0.972 ; 
        RECT 2.34 0.756 2.412 0.972 ; 
        RECT 0.808 0.756 2.412 0.828 ; 
        RECT 0.936 0.252 1.008 0.828 ; 
        RECT 0.808 0.252 1.008 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.104 0.108 2.652 0.18 ; 
      RECT 1.456 0.324 2.432 0.396 ; 
      RECT 0.16 0.9 2.216 0.972 ; 
      RECT 0.376 0.108 1.788 0.18 ; 
  END 
END AOI31xp67_ASAP7_75t_R 


MACRO AOI321xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI321xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.136 0.576 0.656 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.136 0.144 0.944 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.756 1.656 0.828 ; 
        RECT 1.584 0.108 1.656 0.828 ; 
        RECT 0.792 0.108 1.656 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.024 0.9 1.584 0.972 ; 
      RECT 0.376 0.756 0.92 0.828 ; 
  END 
END AOI321xp33_ASAP7_75t_R 


MACRO AOI322xp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI322xp5_ASAP7_75t_R 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.66 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.136 0.36 0.656 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.656 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.66 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.944 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.456 0.756 1.872 0.828 ; 
        RECT 1.8 0.108 1.872 0.828 ; 
        RECT 0.588 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.808 0.9 1.8 0.972 ; 
      RECT 0.156 0.756 1.136 0.828 ; 
  END 
END AOI322xp5_ASAP7_75t_R 


MACRO AOI32xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI32xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.232 0.972 ; 
        RECT 0.072 0.252 0.232 0.324 ; 
        RECT 0.072 0.252 0.144 0.972 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.416 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.416 0.252 0.576 0.324 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.756 0.888 0.828 ; 
        RECT 0.72 0.28 0.792 0.828 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.656 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.756 1.44 0.828 ; 
        RECT 1.368 0.108 1.44 0.828 ; 
        RECT 0.16 0.108 1.44 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.9 1.352 0.972 ; 
  END 
END AOI32xp33_ASAP7_75t_R 


MACRO AOI331xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI331xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.136 0.576 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.136 0.36 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.656 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.656 ; 
    END 
  END C1 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.944 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.668 0.9 1.872 0.972 ; 
        RECT 1.8 0.108 1.872 0.972 ; 
        RECT 0.804 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.016 0.756 1.572 0.828 ; 
      RECT 0.368 0.9 1.356 0.972 ; 
  END 
END AOI331xp33_ASAP7_75t_R 


MACRO AOI332xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI332xp33_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.136 0.576 0.656 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.136 0.36 0.656 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.656 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.28 1.872 0.656 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.656 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.668 0.756 2.088 0.828 ; 
        RECT 2.016 0.108 2.088 0.828 ; 
        RECT 0.804 0.108 2.088 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.016 0.9 2.008 0.972 ; 
      RECT 0.368 0.756 1.356 0.828 ; 
  END 
END AOI332xp33_ASAP7_75t_R 


MACRO AOI333xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI333xp33_ASAP7_75t_R 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.28 2.088 0.656 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.28 1.872 0.656 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.656 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.656 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.136 0.576 0.656 ; 
    END 
  END C2 
  PIN C3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.136 0.36 0.656 ; 
    END 
  END C3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.652 0.756 2.304 0.828 ; 
        RECT 2.232 0.108 2.304 0.828 ; 
        RECT 0.804 0.108 2.304 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.016 0.9 2.06 0.972 ; 
      RECT 0.376 0.756 1.36 0.828 ; 
  END 
END AOI333xp33_ASAP7_75t_R 


MACRO AOI33xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN AOI33xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.136 0.36 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.136 0.576 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.656 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.656 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END B3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.756 1.656 0.828 ; 
        RECT 1.584 0.108 1.656 0.828 ; 
        RECT 0.804 0.108 1.656 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.9 1.352 0.972 ; 
  END 
END AOI33xp33_ASAP7_75t_R 


MACRO ASYNC_DFFHx1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ASYNC_DFFHx1_ASAP7_75t_R 0 0 ; 
  SIZE 5.616 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.728 0.468 0.944 ; 
        RECT 0.288 0.28 0.468 0.352 ; 
        RECT 0.396 0.136 0.468 0.352 ; 
        RECT 0.288 0.728 0.468 0.8 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.504 1.16 0.576 ; 
        RECT 0.936 0.9 1.084 0.972 ; 
        RECT 0.936 0.108 1.084 0.18 ; 
        RECT 0.936 0.108 1.008 0.972 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.344 0.9 5.544 0.972 ; 
        RECT 5.472 0.108 5.544 0.972 ; 
        RECT 5.344 0.108 5.544 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 5.616 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.616 0.036 ; 
    END 
  END VSS 
  PIN RESET 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 2.528 0.432 4.268 0.504 ; 
      LAYER M1 ; 
        RECT 4.176 0.412 4.248 0.672 ; 
        RECT 2.448 0.72 2.672 0.792 ; 
        RECT 2.448 0.432 2.648 0.504 ; 
        RECT 2.448 0.432 2.52 0.792 ; 
      LAYER V1 ; 
        RECT 2.548 0.432 2.62 0.504 ; 
        RECT 4.176 0.432 4.248 0.504 ; 
    END 
  END RESET 
  PIN SET 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 3.132 0.288 4.268 0.36 ; 
      LAYER M1 ; 
        RECT 3.096 0.288 3.244 0.36 ; 
        RECT 3.096 0.288 3.168 0.692 ; 
      LAYER V1 ; 
        RECT 3.152 0.288 3.224 0.36 ; 
    END 
  END SET 
  OBS 
    LAYER M1 ; 
      RECT 3.852 0.864 4.032 0.936 ; 
      RECT 3.852 0.144 3.924 0.936 ; 
      RECT 3.672 0.12 3.744 0.868 ; 
      RECT 3.432 0.12 3.744 0.192 ; 
      RECT 2.232 0.864 3.08 0.936 ; 
      RECT 2.772 0.232 2.844 0.936 ; 
      RECT 2.232 0.656 2.304 0.936 ; 
      RECT 1.672 0.9 2.016 0.972 ; 
      RECT 1.944 0.288 2.016 0.972 ; 
      RECT 1.944 0.288 2.188 0.36 ; 
      RECT 0.592 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.592 0.108 0.792 0.18 ; 
      RECT 0.072 0.9 0.272 0.972 ; 
      RECT 0.072 0.108 0.144 0.972 ; 
      RECT 0.072 0.576 0.188 0.648 ; 
      RECT 0.072 0.108 0.272 0.18 ; 
      RECT 5.256 0.36 5.328 0.668 ; 
      RECT 4.68 0.144 4.808 0.216 ; 
      RECT 4.392 0.412 4.464 0.672 ; 
      RECT 3.528 0.388 3.6 0.812 ; 
      RECT 3.316 0.396 3.388 0.668 ; 
      RECT 3.112 0.144 3.276 0.216 ; 
      RECT 2.916 0.268 2.988 0.532 ; 
      RECT 1.66 0.108 2.432 0.18 ; 
      RECT 1.8 0.476 1.872 0.668 ; 
      RECT 1.584 0.48 1.656 0.812 ; 
      RECT 1.476 0.216 1.548 0.404 ; 
      RECT 1.368 0.48 1.44 0.668 ; 
      RECT 0.568 0.424 0.64 0.668 ; 
    LAYER M2 ; 
      RECT 3.652 0.576 5.348 0.648 ; 
      RECT 3.132 0.144 4.792 0.216 ; 
      RECT 2.964 0.864 4.032 0.936 ; 
      RECT 0.7 0.72 3.704 0.792 ; 
      RECT 0.076 0.576 3.408 0.648 ; 
      RECT 1.456 0.288 3.008 0.36 ; 
    LAYER V1 ; 
      RECT 5.256 0.576 5.328 0.648 ; 
      RECT 4.7 0.144 4.772 0.216 ; 
      RECT 4.392 0.576 4.464 0.648 ; 
      RECT 3.94 0.864 4.012 0.936 ; 
      RECT 3.672 0.576 3.744 0.648 ; 
      RECT 3.528 0.72 3.6 0.792 ; 
      RECT 3.316 0.576 3.388 0.648 ; 
      RECT 3.152 0.144 3.224 0.216 ; 
      RECT 2.984 0.864 3.056 0.936 ; 
      RECT 2.916 0.288 2.988 0.36 ; 
      RECT 2.048 0.288 2.12 0.36 ; 
      RECT 1.8 0.576 1.872 0.648 ; 
      RECT 1.584 0.72 1.656 0.792 ; 
      RECT 1.476 0.288 1.548 0.36 ; 
      RECT 1.368 0.576 1.44 0.648 ; 
      RECT 0.72 0.72 0.792 0.792 ; 
      RECT 0.568 0.576 0.64 0.648 ; 
      RECT 0.096 0.576 0.168 0.648 ; 
  END 
END ASYNC_DFFHx1_ASAP7_75t_R 


MACRO BUFx10_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx10_ASAP7_75t_R 0 0 ; 
  SIZE 3.024 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.024 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.796 0.9 2.952 0.972 ; 
        RECT 2.88 0.108 2.952 0.972 ; 
        RECT 0.796 0.108 2.952 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.364 0.9 0.576 0.972 ; 
      RECT 0.504 0.108 0.576 0.972 ; 
      RECT 0.504 0.504 2.756 0.576 ; 
      RECT 0.364 0.108 0.576 0.18 ; 
  END 
END BUFx10_ASAP7_75t_R 


MACRO BUFx12_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx12_ASAP7_75t_R 0 0 ; 
  SIZE 3.456 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.456 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.456 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.796 0.9 3.384 0.972 ; 
        RECT 3.312 0.108 3.384 0.972 ; 
        RECT 0.796 0.108 3.384 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.9 0.576 0.972 ; 
      RECT 0.504 0.108 0.576 0.972 ; 
      RECT 0.504 0.504 3.2 0.576 ; 
      RECT 0.376 0.108 0.576 0.18 ; 
  END 
END BUFx12_ASAP7_75t_R 


MACRO BUFx12f_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx12f_ASAP7_75t_R 0 0 ; 
  SIZE 3.888 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.296 0.576 ; 
        RECT 0.072 0.136 0.144 0.944 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.888 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.888 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.9 3.816 0.972 ; 
        RECT 3.744 0.108 3.816 0.972 ; 
        RECT 1.24 0.108 3.816 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.9 1.116 0.972 ; 
      RECT 1.044 0.108 1.116 0.972 ; 
      RECT 1.044 0.504 1.244 0.576 ; 
      RECT 0.376 0.108 1.116 0.18 ; 
  END 
END BUFx12f_ASAP7_75t_R 


MACRO BUFx16f_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx16f_ASAP7_75t_R 0 0 ; 
  SIZE 4.752 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.24 0.972 ; 
        RECT 0.072 0.108 0.24 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.752 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.752 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.9 4.68 0.972 ; 
        RECT 4.608 0.108 4.68 0.972 ; 
        RECT 1.24 0.108 4.68 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.9 1.008 0.972 ; 
      RECT 0.936 0.108 1.008 0.972 ; 
      RECT 0.936 0.504 4.496 0.576 ; 
      RECT 0.376 0.108 1.008 0.18 ; 
  END 
END BUFx16f_ASAP7_75t_R 


MACRO BUFx24_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx24_ASAP7_75t_R 0 0 ; 
  SIZE 6.48 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 6.48 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.48 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.9 6.408 0.972 ; 
        RECT 6.336 0.108 6.408 0.972 ; 
        RECT 1.24 0.108 6.408 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.9 1.008 0.972 ; 
      RECT 0.936 0.108 1.008 0.972 ; 
      RECT 0.936 0.504 6.212 0.576 ; 
      RECT 0.376 0.108 1.008 0.18 ; 
  END 
END BUFx24_ASAP7_75t_R 


MACRO BUFx2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx2_ASAP7_75t_R 0 0 ; 
  SIZE 1.08 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.292 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.828 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.08 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.58 0.9 1.008 0.972 ; 
        RECT 0.936 0.108 1.008 0.972 ; 
        RECT 0.58 0.108 1.008 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.48 0.972 ; 
      RECT 0.408 0.108 0.48 0.972 ; 
      RECT 0.408 0.504 0.812 0.576 ; 
      RECT 0.16 0.108 0.48 0.18 ; 
  END 
END BUFx2_ASAP7_75t_R 


MACRO BUFx3_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx3_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.292 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.828 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.58 0.9 1.224 0.972 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
        RECT 0.58 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.48 0.972 ; 
      RECT 0.408 0.108 0.48 0.972 ; 
      RECT 0.408 0.504 1.04 0.576 ; 
      RECT 0.16 0.108 0.48 0.18 ; 
  END 
END BUFx3_ASAP7_75t_R 


MACRO BUFx4_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx4_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.292 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.828 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.58 0.9 1.428 0.972 ; 
        RECT 1.356 0.108 1.428 0.972 ; 
        RECT 0.58 0.108 1.428 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.48 0.972 ; 
      RECT 0.408 0.108 0.48 0.972 ; 
      RECT 0.408 0.504 1.256 0.576 ; 
      RECT 0.16 0.108 0.48 0.18 ; 
  END 
END BUFx4_ASAP7_75t_R 


MACRO BUFx4f_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx4f_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.392 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.796 0.9 1.656 0.972 ; 
        RECT 1.584 0.108 1.656 0.972 ; 
        RECT 0.796 0.108 1.656 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.364 0.9 0.576 0.972 ; 
      RECT 0.504 0.108 0.576 0.972 ; 
      RECT 0.504 0.504 1.468 0.576 ; 
      RECT 0.364 0.108 0.576 0.18 ; 
  END 
END BUFx4f_ASAP7_75t_R 


MACRO BUFx5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx5_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.292 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.828 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.58 0.9 1.656 0.972 ; 
        RECT 1.584 0.108 1.656 0.972 ; 
        RECT 0.58 0.108 1.656 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.48 0.972 ; 
      RECT 0.408 0.108 0.48 0.972 ; 
      RECT 0.408 0.504 1.472 0.576 ; 
      RECT 0.16 0.108 0.48 0.18 ; 
  END 
END BUFx5_ASAP7_75t_R 


MACRO BUFx6f_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx6f_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.336 0.576 ; 
        RECT 0.072 0.136 0.144 0.944 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.9 2.088 0.972 ; 
        RECT 2.016 0.108 2.088 0.972 ; 
        RECT 0.808 0.108 2.088 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.9 0.576 0.972 ; 
      RECT 0.504 0.108 0.576 0.972 ; 
      RECT 0.504 0.504 1.892 0.576 ; 
      RECT 0.376 0.108 0.576 0.18 ; 
  END 
END BUFx6f_ASAP7_75t_R 


MACRO BUFx8_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN BUFx8_ASAP7_75t_R 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.392 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.592 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.9 2.52 0.972 ; 
        RECT 2.448 0.108 2.52 0.972 ; 
        RECT 0.808 0.108 2.52 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.364 0.9 0.576 0.972 ; 
      RECT 0.504 0.108 0.576 0.972 ; 
      RECT 0.504 0.504 2.324 0.576 ; 
      RECT 0.364 0.108 0.576 0.18 ; 
  END 
END BUFx8_ASAP7_75t_R 


MACRO CKINVDCx10_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx10_ASAP7_75t_R 0 0 ; 
  SIZE 5.184 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.352 0.504 4.68 0.576 ; 
        RECT 4.48 0.108 4.552 0.576 ; 
        RECT 0.2 0.108 4.552 0.18 ; 
        RECT 3.056 0.504 3.256 0.576 ; 
        RECT 3.184 0.108 3.256 0.576 ; 
        RECT 1.496 0.504 1.696 0.576 ; 
        RECT 1.496 0.108 1.568 0.576 ; 
        RECT 0.2 0.504 0.4 0.576 ; 
        RECT 0.2 0.108 0.272 0.576 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 5.184 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.184 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 4.896 0.972 ; 
        RECT 4.824 0.252 4.896 0.972 ; 
        RECT 4.696 0.252 4.896 0.324 ; 
        RECT 4.176 0.252 4.376 0.324 ; 
        RECT 4.176 0.252 4.248 0.972 ; 
        RECT 2.88 0.252 3.08 0.324 ; 
        RECT 2.88 0.252 2.952 0.972 ; 
        RECT 1.8 0.252 1.872 0.972 ; 
        RECT 1.672 0.252 1.872 0.324 ; 
        RECT 0.504 0.252 0.576 0.972 ; 
        RECT 0.376 0.252 0.576 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 3.744 0.504 3.968 0.576 ; 
      RECT 3.744 0.36 3.816 0.576 ; 
      RECT 3.4 0.36 4.008 0.432 ; 
      RECT 3.324 0.648 3.944 0.72 ; 
      RECT 3.528 0.504 3.6 0.72 ; 
      RECT 3.368 0.504 3.6 0.576 ; 
      RECT 2.104 0.648 2.724 0.72 ; 
      RECT 2.448 0.504 2.52 0.72 ; 
      RECT 2.448 0.504 2.68 0.576 ; 
      RECT 2.08 0.504 2.304 0.576 ; 
      RECT 2.232 0.36 2.304 0.576 ; 
      RECT 2.04 0.36 2.648 0.432 ; 
      RECT 0.808 0.648 1.428 0.72 ; 
      RECT 1.152 0.504 1.224 0.72 ; 
      RECT 1.152 0.504 1.384 0.576 ; 
      RECT 0.784 0.504 1.008 0.576 ; 
      RECT 0.936 0.36 1.008 0.576 ; 
      RECT 0.744 0.36 1.352 0.432 ; 
  END 
END CKINVDCx10_ASAP7_75t_R 


MACRO CKINVDCx11_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx11_ASAP7_75t_R 0 0 ; 
  SIZE 5.616 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.216 0.504 5.416 0.576 ; 
        RECT 5.344 0.108 5.416 0.576 ; 
        RECT 0.2 0.108 5.416 0.18 ; 
        RECT 3.488 0.504 3.856 0.576 ; 
        RECT 3.636 0.108 3.708 0.576 ; 
        RECT 1.756 0.504 2.124 0.576 ; 
        RECT 1.904 0.108 1.976 0.576 ; 
        RECT 0.2 0.504 0.4 0.576 ; 
        RECT 0.2 0.108 0.272 0.576 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 5.616 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.616 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 5.24 0.972 ; 
        RECT 5.04 0.252 5.24 0.324 ; 
        RECT 5.04 0.252 5.112 0.972 ; 
        RECT 3.96 0.252 4.032 0.972 ; 
        RECT 3.832 0.252 4.032 0.324 ; 
        RECT 3.312 0.252 3.512 0.324 ; 
        RECT 3.312 0.252 3.384 0.972 ; 
        RECT 2.232 0.252 2.304 0.972 ; 
        RECT 2.104 0.252 2.304 0.324 ; 
        RECT 1.584 0.252 1.784 0.324 ; 
        RECT 1.584 0.252 1.656 0.972 ; 
        RECT 0.504 0.252 0.576 0.972 ; 
        RECT 0.376 0.252 0.576 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.504 4.832 0.576 ; 
      RECT 4.608 0.36 4.68 0.576 ; 
      RECT 4.264 0.36 4.872 0.432 ; 
      RECT 4.188 0.648 4.808 0.72 ; 
      RECT 4.392 0.504 4.464 0.72 ; 
      RECT 4.232 0.504 4.464 0.576 ; 
      RECT 2.536 0.648 3.156 0.72 ; 
      RECT 2.88 0.504 2.952 0.72 ; 
      RECT 2.88 0.504 3.112 0.576 ; 
      RECT 2.512 0.504 2.736 0.576 ; 
      RECT 2.664 0.36 2.736 0.576 ; 
      RECT 2.472 0.36 3.08 0.432 ; 
      RECT 0.808 0.648 1.428 0.72 ; 
      RECT 1.152 0.504 1.224 0.72 ; 
      RECT 1.152 0.504 1.384 0.576 ; 
      RECT 0.784 0.504 1.008 0.576 ; 
      RECT 0.936 0.36 1.008 0.576 ; 
      RECT 0.744 0.36 1.352 0.432 ; 
  END 
END CKINVDCx11_ASAP7_75t_R 


MACRO CKINVDCx12_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx12_ASAP7_75t_R 0 0 ; 
  SIZE 5.616 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.216 0.504 5.416 0.576 ; 
        RECT 5.344 0.108 5.416 0.576 ; 
        RECT 0.2 0.108 5.416 0.18 ; 
        RECT 3.488 0.504 3.856 0.576 ; 
        RECT 3.636 0.108 3.708 0.576 ; 
        RECT 1.756 0.504 2.124 0.576 ; 
        RECT 1.904 0.108 1.976 0.576 ; 
        RECT 0.2 0.504 0.4 0.576 ; 
        RECT 0.2 0.108 0.272 0.576 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 5.616 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.616 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 5.24 0.972 ; 
        RECT 5.04 0.252 5.24 0.324 ; 
        RECT 5.04 0.252 5.112 0.972 ; 
        RECT 3.96 0.252 4.032 0.972 ; 
        RECT 3.832 0.252 4.032 0.324 ; 
        RECT 3.312 0.252 3.512 0.324 ; 
        RECT 3.312 0.252 3.384 0.972 ; 
        RECT 2.232 0.252 2.304 0.972 ; 
        RECT 2.104 0.252 2.304 0.324 ; 
        RECT 1.584 0.252 1.784 0.324 ; 
        RECT 1.584 0.252 1.656 0.972 ; 
        RECT 0.504 0.252 0.576 0.972 ; 
        RECT 0.376 0.252 0.576 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.504 4.832 0.576 ; 
      RECT 4.608 0.36 4.68 0.576 ; 
      RECT 4.264 0.36 4.872 0.432 ; 
      RECT 4.188 0.648 4.808 0.72 ; 
      RECT 4.392 0.504 4.464 0.72 ; 
      RECT 4.232 0.504 4.464 0.576 ; 
      RECT 2.536 0.648 3.156 0.72 ; 
      RECT 2.88 0.504 2.952 0.72 ; 
      RECT 2.88 0.504 3.112 0.576 ; 
      RECT 2.512 0.504 2.736 0.576 ; 
      RECT 2.664 0.36 2.736 0.576 ; 
      RECT 2.472 0.36 3.08 0.432 ; 
      RECT 0.808 0.648 1.428 0.72 ; 
      RECT 1.152 0.504 1.224 0.72 ; 
      RECT 1.152 0.504 1.384 0.576 ; 
      RECT 0.784 0.504 1.008 0.576 ; 
      RECT 0.936 0.36 1.008 0.576 ; 
      RECT 0.744 0.36 1.352 0.432 ; 
  END 
END CKINVDCx12_ASAP7_75t_R 


MACRO CKINVDCx14_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx14_ASAP7_75t_R 0 0 ; 
  SIZE 6.048 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.216 0.504 5.588 0.576 ; 
        RECT 5.344 0.108 5.416 0.576 ; 
        RECT 0.2 0.108 5.416 0.18 ; 
        RECT 3.488 0.504 3.856 0.576 ; 
        RECT 3.636 0.108 3.708 0.576 ; 
        RECT 1.756 0.504 2.124 0.576 ; 
        RECT 1.904 0.108 1.976 0.576 ; 
        RECT 0.2 0.504 0.4 0.576 ; 
        RECT 0.2 0.108 0.272 0.576 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 6.048 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.048 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 5.76 0.972 ; 
        RECT 5.688 0.252 5.76 0.972 ; 
        RECT 5.56 0.252 5.76 0.324 ; 
        RECT 5.04 0.252 5.24 0.324 ; 
        RECT 5.04 0.252 5.112 0.972 ; 
        RECT 3.96 0.252 4.032 0.972 ; 
        RECT 3.832 0.252 4.032 0.324 ; 
        RECT 3.312 0.252 3.512 0.324 ; 
        RECT 3.312 0.252 3.384 0.972 ; 
        RECT 2.232 0.252 2.304 0.972 ; 
        RECT 2.104 0.252 2.304 0.324 ; 
        RECT 1.584 0.252 1.784 0.324 ; 
        RECT 1.584 0.252 1.656 0.972 ; 
        RECT 0.504 0.252 0.576 0.972 ; 
        RECT 0.376 0.252 0.576 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.504 4.832 0.576 ; 
      RECT 4.608 0.36 4.68 0.576 ; 
      RECT 4.264 0.36 4.872 0.432 ; 
      RECT 4.188 0.648 4.808 0.72 ; 
      RECT 4.392 0.504 4.464 0.72 ; 
      RECT 4.232 0.504 4.464 0.576 ; 
      RECT 2.536 0.648 3.156 0.72 ; 
      RECT 2.88 0.504 2.952 0.72 ; 
      RECT 2.88 0.504 3.112 0.576 ; 
      RECT 2.512 0.504 2.736 0.576 ; 
      RECT 2.664 0.36 2.736 0.576 ; 
      RECT 2.472 0.36 3.08 0.432 ; 
      RECT 0.808 0.648 1.428 0.72 ; 
      RECT 1.152 0.504 1.224 0.72 ; 
      RECT 1.152 0.504 1.384 0.576 ; 
      RECT 0.784 0.504 1.008 0.576 ; 
      RECT 0.936 0.36 1.008 0.576 ; 
      RECT 0.744 0.36 1.352 0.432 ; 
  END 
END CKINVDCx14_ASAP7_75t_R 


MACRO CKINVDCx16_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx16_ASAP7_75t_R 0 0 ; 
  SIZE 6.48 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.648 0.504 6.02 0.576 ; 
        RECT 5.776 0.108 5.848 0.576 ; 
        RECT 0.632 0.108 5.848 0.18 ; 
        RECT 3.92 0.504 4.288 0.576 ; 
        RECT 4.068 0.108 4.14 0.576 ; 
        RECT 2.188 0.504 2.556 0.576 ; 
        RECT 2.336 0.108 2.408 0.576 ; 
        RECT 0.504 0.504 0.832 0.576 ; 
        RECT 0.632 0.108 0.704 0.576 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 6.48 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.48 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.9 6.192 0.972 ; 
        RECT 6.12 0.252 6.192 0.972 ; 
        RECT 5.992 0.252 6.192 0.324 ; 
        RECT 5.472 0.252 5.672 0.324 ; 
        RECT 5.472 0.252 5.544 0.972 ; 
        RECT 4.392 0.252 4.464 0.972 ; 
        RECT 4.264 0.252 4.464 0.324 ; 
        RECT 3.744 0.252 3.944 0.324 ; 
        RECT 3.744 0.252 3.816 0.972 ; 
        RECT 2.664 0.252 2.736 0.972 ; 
        RECT 2.536 0.252 2.736 0.324 ; 
        RECT 2.016 0.252 2.216 0.324 ; 
        RECT 2.016 0.252 2.088 0.972 ; 
        RECT 0.936 0.252 1.008 0.972 ; 
        RECT 0.808 0.252 1.008 0.324 ; 
        RECT 0.288 0.252 0.488 0.324 ; 
        RECT 0.288 0.252 0.36 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 5.04 0.504 5.264 0.576 ; 
      RECT 5.04 0.36 5.112 0.576 ; 
      RECT 4.696 0.36 5.304 0.432 ; 
      RECT 4.62 0.648 5.24 0.72 ; 
      RECT 4.824 0.504 4.896 0.72 ; 
      RECT 4.664 0.504 4.896 0.576 ; 
      RECT 2.968 0.648 3.588 0.72 ; 
      RECT 3.312 0.504 3.384 0.72 ; 
      RECT 3.312 0.504 3.544 0.576 ; 
      RECT 2.944 0.504 3.168 0.576 ; 
      RECT 3.096 0.36 3.168 0.576 ; 
      RECT 2.904 0.36 3.512 0.432 ; 
      RECT 1.24 0.648 1.86 0.72 ; 
      RECT 1.584 0.504 1.656 0.72 ; 
      RECT 1.584 0.504 1.816 0.576 ; 
      RECT 1.216 0.504 1.44 0.576 ; 
      RECT 1.368 0.36 1.44 0.576 ; 
      RECT 1.176 0.36 1.784 0.432 ; 
  END 
END CKINVDCx16_ASAP7_75t_R 


MACRO CKINVDCx20_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx20_ASAP7_75t_R 0 0 ; 
  SIZE 8.208 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 7.376 0.504 7.748 0.576 ; 
        RECT 7.504 0.108 7.576 0.576 ; 
        RECT 0.632 0.108 7.576 0.18 ; 
        RECT 5.648 0.504 6.02 0.576 ; 
        RECT 5.776 0.108 5.848 0.576 ; 
        RECT 3.92 0.504 4.288 0.576 ; 
        RECT 4.068 0.108 4.14 0.576 ; 
        RECT 2.188 0.504 2.556 0.576 ; 
        RECT 2.336 0.108 2.408 0.576 ; 
        RECT 0.504 0.504 0.832 0.576 ; 
        RECT 0.632 0.108 0.704 0.576 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 8.208 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 8.208 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.9 7.92 0.972 ; 
        RECT 7.848 0.252 7.92 0.972 ; 
        RECT 7.72 0.252 7.92 0.324 ; 
        RECT 7.2 0.252 7.4 0.324 ; 
        RECT 7.2 0.252 7.272 0.972 ; 
        RECT 6.12 0.252 6.192 0.972 ; 
        RECT 5.992 0.252 6.192 0.324 ; 
        RECT 5.472 0.252 5.672 0.324 ; 
        RECT 5.472 0.252 5.544 0.972 ; 
        RECT 4.392 0.252 4.464 0.972 ; 
        RECT 4.264 0.252 4.464 0.324 ; 
        RECT 3.744 0.252 3.944 0.324 ; 
        RECT 3.744 0.252 3.816 0.972 ; 
        RECT 2.664 0.252 2.736 0.972 ; 
        RECT 2.536 0.252 2.736 0.324 ; 
        RECT 2.016 0.252 2.216 0.324 ; 
        RECT 2.016 0.252 2.088 0.972 ; 
        RECT 0.936 0.252 1.008 0.972 ; 
        RECT 0.808 0.252 1.008 0.324 ; 
        RECT 0.288 0.252 0.488 0.324 ; 
        RECT 0.288 0.252 0.36 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 6.768 0.504 6.992 0.576 ; 
      RECT 6.768 0.36 6.84 0.576 ; 
      RECT 6.424 0.36 7.032 0.432 ; 
      RECT 6.348 0.648 6.968 0.72 ; 
      RECT 6.552 0.504 6.624 0.72 ; 
      RECT 6.392 0.504 6.624 0.576 ; 
      RECT 5.04 0.504 5.264 0.576 ; 
      RECT 5.04 0.36 5.112 0.576 ; 
      RECT 4.696 0.36 5.304 0.432 ; 
      RECT 4.62 0.648 5.24 0.72 ; 
      RECT 4.824 0.504 4.896 0.72 ; 
      RECT 4.664 0.504 4.896 0.576 ; 
      RECT 2.968 0.648 3.588 0.72 ; 
      RECT 3.312 0.504 3.384 0.72 ; 
      RECT 3.312 0.504 3.544 0.576 ; 
      RECT 2.944 0.504 3.168 0.576 ; 
      RECT 3.096 0.36 3.168 0.576 ; 
      RECT 2.904 0.36 3.512 0.432 ; 
      RECT 1.24 0.648 1.86 0.72 ; 
      RECT 1.584 0.504 1.656 0.72 ; 
      RECT 1.584 0.504 1.816 0.576 ; 
      RECT 1.216 0.504 1.44 0.576 ; 
      RECT 1.368 0.36 1.44 0.576 ; 
      RECT 1.176 0.36 1.784 0.432 ; 
  END 
END CKINVDCx20_ASAP7_75t_R 


MACRO CKINVDCx5p33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx5p33_ASAP7_75t_R 0 0 ; 
  SIZE 4.752 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.352 0.504 4.552 0.576 ; 
        RECT 4.48 0.108 4.552 0.576 ; 
        RECT 0.2 0.108 4.552 0.18 ; 
        RECT 3.056 0.504 3.256 0.576 ; 
        RECT 3.184 0.108 3.256 0.576 ; 
        RECT 1.496 0.504 1.696 0.576 ; 
        RECT 1.496 0.108 1.568 0.576 ; 
        RECT 0.2 0.504 0.4 0.576 ; 
        RECT 0.2 0.108 0.272 0.576 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.752 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.752 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 4.376 0.972 ; 
        RECT 4.176 0.252 4.376 0.324 ; 
        RECT 4.176 0.252 4.248 0.972 ; 
        RECT 2.88 0.252 3.08 0.324 ; 
        RECT 2.88 0.252 2.952 0.972 ; 
        RECT 1.8 0.252 1.872 0.972 ; 
        RECT 1.672 0.252 1.872 0.324 ; 
        RECT 0.504 0.252 0.576 0.972 ; 
        RECT 0.376 0.252 0.576 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 3.744 0.504 3.968 0.576 ; 
      RECT 3.744 0.36 3.816 0.576 ; 
      RECT 3.4 0.36 4.008 0.432 ; 
      RECT 3.324 0.648 3.944 0.72 ; 
      RECT 3.528 0.504 3.6 0.72 ; 
      RECT 3.368 0.504 3.6 0.576 ; 
      RECT 2.104 0.648 2.724 0.72 ; 
      RECT 2.448 0.504 2.52 0.72 ; 
      RECT 2.448 0.504 2.68 0.576 ; 
      RECT 2.08 0.504 2.304 0.576 ; 
      RECT 2.232 0.36 2.304 0.576 ; 
      RECT 2.04 0.36 2.648 0.432 ; 
      RECT 0.808 0.648 1.428 0.72 ; 
      RECT 1.152 0.504 1.224 0.72 ; 
      RECT 1.152 0.504 1.384 0.576 ; 
      RECT 0.784 0.504 1.008 0.576 ; 
      RECT 0.936 0.36 1.008 0.576 ; 
      RECT 0.744 0.36 1.352 0.432 ; 
  END 
END CKINVDCx5p33_ASAP7_75t_R 


MACRO CKINVDCx6p67_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx6p67_ASAP7_75t_R 0 0 ; 
  SIZE 5.184 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.352 0.504 4.68 0.576 ; 
        RECT 4.48 0.108 4.552 0.576 ; 
        RECT 0.2 0.108 4.552 0.18 ; 
        RECT 3.056 0.504 3.256 0.576 ; 
        RECT 3.184 0.108 3.256 0.576 ; 
        RECT 1.496 0.504 1.696 0.576 ; 
        RECT 1.496 0.108 1.568 0.576 ; 
        RECT 0.2 0.504 0.4 0.576 ; 
        RECT 0.2 0.108 0.272 0.576 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 5.184 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.184 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 4.896 0.972 ; 
        RECT 4.824 0.252 4.896 0.972 ; 
        RECT 4.696 0.252 4.896 0.324 ; 
        RECT 4.176 0.252 4.376 0.324 ; 
        RECT 4.176 0.252 4.248 0.972 ; 
        RECT 2.88 0.252 3.08 0.324 ; 
        RECT 2.88 0.252 2.952 0.972 ; 
        RECT 1.8 0.252 1.872 0.972 ; 
        RECT 1.672 0.252 1.872 0.324 ; 
        RECT 0.504 0.252 0.576 0.972 ; 
        RECT 0.376 0.252 0.576 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 3.744 0.504 3.968 0.576 ; 
      RECT 3.744 0.36 3.816 0.576 ; 
      RECT 3.4 0.36 4.008 0.432 ; 
      RECT 3.324 0.648 3.944 0.72 ; 
      RECT 3.528 0.504 3.6 0.72 ; 
      RECT 3.368 0.504 3.6 0.576 ; 
      RECT 2.104 0.648 2.724 0.72 ; 
      RECT 2.448 0.504 2.52 0.72 ; 
      RECT 2.448 0.504 2.68 0.576 ; 
      RECT 2.08 0.504 2.304 0.576 ; 
      RECT 2.232 0.36 2.304 0.576 ; 
      RECT 2.04 0.36 2.648 0.432 ; 
      RECT 0.808 0.648 1.428 0.72 ; 
      RECT 1.152 0.504 1.224 0.72 ; 
      RECT 1.152 0.504 1.384 0.576 ; 
      RECT 0.784 0.504 1.008 0.576 ; 
      RECT 0.936 0.36 1.008 0.576 ; 
      RECT 0.744 0.36 1.352 0.432 ; 
  END 
END CKINVDCx6p67_ASAP7_75t_R 


MACRO CKINVDCx8_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx8_ASAP7_75t_R 0 0 ; 
  SIZE 4.752 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.352 0.504 4.552 0.576 ; 
        RECT 4.48 0.108 4.552 0.576 ; 
        RECT 0.2 0.108 4.552 0.18 ; 
        RECT 3.056 0.504 3.256 0.576 ; 
        RECT 3.184 0.108 3.256 0.576 ; 
        RECT 1.496 0.504 1.696 0.576 ; 
        RECT 1.496 0.108 1.568 0.576 ; 
        RECT 0.2 0.504 0.4 0.576 ; 
        RECT 0.2 0.108 0.272 0.576 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.752 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.752 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 4.376 0.972 ; 
        RECT 4.176 0.252 4.376 0.324 ; 
        RECT 4.176 0.252 4.248 0.972 ; 
        RECT 2.88 0.252 3.08 0.324 ; 
        RECT 2.88 0.252 2.952 0.972 ; 
        RECT 1.8 0.252 1.872 0.972 ; 
        RECT 1.672 0.252 1.872 0.324 ; 
        RECT 0.504 0.252 0.576 0.972 ; 
        RECT 0.376 0.252 0.576 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 3.744 0.504 3.968 0.576 ; 
      RECT 3.744 0.36 3.816 0.576 ; 
      RECT 3.4 0.36 4.008 0.432 ; 
      RECT 3.324 0.648 3.944 0.72 ; 
      RECT 3.528 0.504 3.6 0.72 ; 
      RECT 3.368 0.504 3.6 0.576 ; 
      RECT 2.104 0.648 2.724 0.72 ; 
      RECT 2.448 0.504 2.52 0.72 ; 
      RECT 2.448 0.504 2.68 0.576 ; 
      RECT 2.08 0.504 2.304 0.576 ; 
      RECT 2.232 0.36 2.304 0.576 ; 
      RECT 2.04 0.36 2.648 0.432 ; 
      RECT 0.808 0.648 1.428 0.72 ; 
      RECT 1.152 0.504 1.224 0.72 ; 
      RECT 1.152 0.504 1.384 0.576 ; 
      RECT 0.784 0.504 1.008 0.576 ; 
      RECT 0.936 0.36 1.008 0.576 ; 
      RECT 0.744 0.36 1.352 0.432 ; 
  END 
END CKINVDCx8_ASAP7_75t_R 


MACRO CKINVDCx9p33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN CKINVDCx9p33_ASAP7_75t_R 0 0 ; 
  SIZE 6.048 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.216 0.504 5.588 0.576 ; 
        RECT 5.344 0.108 5.416 0.576 ; 
        RECT 0.2 0.108 5.416 0.18 ; 
        RECT 3.488 0.504 3.856 0.576 ; 
        RECT 3.636 0.108 3.708 0.576 ; 
        RECT 1.756 0.504 2.124 0.576 ; 
        RECT 1.904 0.108 1.976 0.576 ; 
        RECT 0.2 0.504 0.4 0.576 ; 
        RECT 0.2 0.108 0.272 0.576 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 6.048 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.048 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 5.76 0.972 ; 
        RECT 5.688 0.252 5.76 0.972 ; 
        RECT 5.56 0.252 5.76 0.324 ; 
        RECT 5.04 0.252 5.24 0.324 ; 
        RECT 5.04 0.252 5.112 0.972 ; 
        RECT 3.96 0.252 4.032 0.972 ; 
        RECT 3.832 0.252 4.032 0.324 ; 
        RECT 3.312 0.252 3.512 0.324 ; 
        RECT 3.312 0.252 3.384 0.972 ; 
        RECT 2.232 0.252 2.304 0.972 ; 
        RECT 2.104 0.252 2.304 0.324 ; 
        RECT 1.584 0.252 1.784 0.324 ; 
        RECT 1.584 0.252 1.656 0.972 ; 
        RECT 0.504 0.252 0.576 0.972 ; 
        RECT 0.376 0.252 0.576 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.504 4.832 0.576 ; 
      RECT 4.608 0.36 4.68 0.576 ; 
      RECT 4.264 0.36 4.872 0.432 ; 
      RECT 4.188 0.648 4.808 0.72 ; 
      RECT 4.392 0.504 4.464 0.72 ; 
      RECT 4.232 0.504 4.464 0.576 ; 
      RECT 2.536 0.648 3.156 0.72 ; 
      RECT 2.88 0.504 2.952 0.72 ; 
      RECT 2.88 0.504 3.112 0.576 ; 
      RECT 2.512 0.504 2.736 0.576 ; 
      RECT 2.664 0.36 2.736 0.576 ; 
      RECT 2.472 0.36 3.08 0.432 ; 
      RECT 0.808 0.648 1.428 0.72 ; 
      RECT 1.152 0.504 1.224 0.72 ; 
      RECT 1.152 0.504 1.384 0.576 ; 
      RECT 0.784 0.504 1.008 0.576 ; 
      RECT 0.936 0.36 1.008 0.576 ; 
      RECT 0.744 0.36 1.352 0.432 ; 
  END 
END CKINVDCx9p33_ASAP7_75t_R 


MACRO DECAPx10_ASAP7_75t_R 
  CLASS CORE SPACER ; 
  ORIGIN 0 0 ; 
  FOREIGN DECAPx10_ASAP7_75t_R 0 0 ; 
  SIZE 4.752 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.752 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.752 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.232 0.18 2.304 0.6 ; 
      RECT 2.232 0.18 4.592 0.252 ; 
      RECT 0.16 0.828 2.52 0.9 ; 
      RECT 2.448 0.484 2.52 0.9 ; 
  END 
END DECAPx10_ASAP7_75t_R 


MACRO DECAPx1_ASAP7_75t_R 
  CLASS CORE SPACER ; 
  ORIGIN 0 0 ; 
  FOREIGN DECAPx1_ASAP7_75t_R 0 0 ; 
  SIZE 0.864 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.864 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.864 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.828 0.576 0.9 ; 
      RECT 0.504 0.484 0.576 0.9 ; 
      RECT 0.288 0.18 0.36 0.6 ; 
      RECT 0.288 0.18 0.488 0.252 ; 
  END 
END DECAPx1_ASAP7_75t_R 


MACRO DECAPx2_ASAP7_75t_R 
  CLASS CORE SPACER ; 
  ORIGIN 0 0 ; 
  FOREIGN DECAPx2_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 0.504 0.18 0.576 0.6 ; 
      RECT 0.504 0.18 1.136 0.252 ; 
      RECT 0.16 0.828 0.792 0.9 ; 
      RECT 0.72 0.484 0.792 0.9 ; 
  END 
END DECAPx2_ASAP7_75t_R 


MACRO DECAPx2b_ASAP7_75t_R 
  CLASS CORE SPACER ; 
  ORIGIN 0 0 ; 
  FOREIGN DECAPx2b_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.648 0.996 0.72 ; 
      RECT 0.72 0.504 0.792 0.72 ; 
      RECT 0.72 0.504 0.952 0.576 ; 
      RECT 0.352 0.504 0.576 0.576 ; 
      RECT 0.504 0.36 0.576 0.576 ; 
      RECT 0.312 0.36 0.92 0.432 ; 
  END 
END DECAPx2b_ASAP7_75t_R 


MACRO DECAPx4_ASAP7_75t_R 
  CLASS CORE SPACER ; 
  ORIGIN 0 0 ; 
  FOREIGN DECAPx4_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 0.936 0.18 1.008 0.6 ; 
      RECT 0.936 0.18 2 0.252 ; 
      RECT 0.16 0.828 1.224 0.9 ; 
      RECT 1.152 0.484 1.224 0.9 ; 
  END 
END DECAPx4_ASAP7_75t_R 


MACRO DECAPx6_ASAP7_75t_R 
  CLASS CORE SPACER ; 
  ORIGIN 0 0 ; 
  FOREIGN DECAPx6_ASAP7_75t_R 0 0 ; 
  SIZE 3.024 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.024 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 1.368 0.18 1.44 0.6 ; 
      RECT 1.368 0.18 2.864 0.252 ; 
      RECT 0.16 0.828 1.656 0.9 ; 
      RECT 1.584 0.484 1.656 0.9 ; 
  END 
END DECAPx6_ASAP7_75t_R 


MACRO DFFHQNx1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFHQNx1_ASAP7_75t_R 0 0 ; 
  SIZE 4.32 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.656 0.468 0.944 ; 
        RECT 0.288 0.28 0.468 0.424 ; 
        RECT 0.396 0.136 0.468 0.424 ; 
        RECT 0.288 0.656 0.468 0.8 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.504 1.16 0.576 ; 
        RECT 0.936 0.9 1.084 0.972 ; 
        RECT 0.936 0.108 1.084 0.18 ; 
        RECT 0.936 0.108 1.008 0.972 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.048 0.9 4.248 0.972 ; 
        RECT 4.176 0.108 4.248 0.972 ; 
        RECT 4.048 0.108 4.248 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.32 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.32 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 3.4 0.9 3.816 0.972 ; 
      RECT 3.744 0.108 3.816 0.972 ; 
      RECT 3.096 0.108 3.168 0.476 ; 
      RECT 3.096 0.108 3.816 0.18 ; 
      RECT 2.752 0.896 2.952 0.968 ; 
      RECT 2.88 0.108 2.952 0.968 ; 
      RECT 2.88 0.612 3.6 0.684 ; 
      RECT 3.528 0.468 3.6 0.684 ; 
      RECT 3.312 0.468 3.384 0.684 ; 
      RECT 2.536 0.108 2.952 0.18 ; 
      RECT 2.304 0.9 2.52 0.972 ; 
      RECT 2.448 0.324 2.52 0.972 ; 
      RECT 1.984 0.324 2.52 0.396 ; 
      RECT 2.34 0.18 2.412 0.396 ; 
      RECT 1.456 0.9 1.872 0.972 ; 
      RECT 1.8 0.108 1.872 0.972 ; 
      RECT 1.8 0.488 2.304 0.56 ; 
      RECT 1.672 0.108 1.872 0.18 ; 
      RECT 1.26 0.504 1.332 0.812 ; 
      RECT 1.26 0.504 1.468 0.576 ; 
      RECT 0.592 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.592 0.108 0.792 0.18 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.576 0.188 0.648 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 3.96 0.36 4.032 0.668 ; 
      RECT 2.664 0.404 2.736 0.668 ; 
      RECT 2.016 0.66 2.088 0.812 ; 
      RECT 1.584 0.424 1.656 0.668 ; 
      RECT 0.568 0.424 0.64 0.668 ; 
    LAYER M2 ; 
      RECT 3.508 0.576 4.052 0.648 ; 
      RECT 0.076 0.576 2.756 0.648 ; 
      RECT 0.7 0.72 2.108 0.792 ; 
    LAYER V1 ; 
      RECT 3.96 0.576 4.032 0.648 ; 
      RECT 3.528 0.576 3.6 0.648 ; 
      RECT 2.664 0.576 2.736 0.648 ; 
      RECT 2.016 0.72 2.088 0.792 ; 
      RECT 1.584 0.576 1.656 0.648 ; 
      RECT 1.26 0.72 1.332 0.792 ; 
      RECT 0.72 0.72 0.792 0.792 ; 
      RECT 0.568 0.576 0.64 0.648 ; 
      RECT 0.096 0.576 0.168 0.648 ; 
  END 
END DFFHQNx1_ASAP7_75t_R 


MACRO DFFHQNx2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFHQNx2_ASAP7_75t_R 0 0 ; 
  SIZE 4.536 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.656 0.468 0.944 ; 
        RECT 0.288 0.28 0.468 0.424 ; 
        RECT 0.396 0.136 0.468 0.424 ; 
        RECT 0.288 0.656 0.468 0.8 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.504 1.16 0.576 ; 
        RECT 0.936 0.9 1.084 0.972 ; 
        RECT 0.936 0.108 1.084 0.18 ; 
        RECT 0.936 0.108 1.008 0.972 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.048 0.864 4.468 0.936 ; 
        RECT 4.396 0.144 4.468 0.936 ; 
        RECT 4.048 0.144 4.468 0.216 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.536 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.536 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 3.4 0.9 3.816 0.972 ; 
      RECT 3.744 0.108 3.816 0.972 ; 
      RECT 3.096 0.108 3.168 0.476 ; 
      RECT 3.096 0.108 3.816 0.18 ; 
      RECT 2.752 0.896 2.952 0.968 ; 
      RECT 2.88 0.108 2.952 0.968 ; 
      RECT 2.88 0.612 3.6 0.684 ; 
      RECT 3.528 0.468 3.6 0.684 ; 
      RECT 3.312 0.468 3.384 0.684 ; 
      RECT 2.536 0.108 2.952 0.18 ; 
      RECT 2.304 0.9 2.52 0.972 ; 
      RECT 2.448 0.324 2.52 0.972 ; 
      RECT 1.984 0.324 2.52 0.396 ; 
      RECT 2.34 0.18 2.412 0.396 ; 
      RECT 1.456 0.9 1.872 0.972 ; 
      RECT 1.8 0.108 1.872 0.972 ; 
      RECT 1.8 0.488 2.304 0.56 ; 
      RECT 1.672 0.108 1.872 0.18 ; 
      RECT 1.26 0.504 1.332 0.812 ; 
      RECT 1.26 0.504 1.468 0.576 ; 
      RECT 0.592 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.592 0.108 0.792 0.18 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.576 0.188 0.648 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 3.96 0.36 4.032 0.668 ; 
      RECT 2.664 0.404 2.736 0.668 ; 
      RECT 2.016 0.66 2.088 0.812 ; 
      RECT 1.584 0.424 1.656 0.668 ; 
      RECT 0.568 0.424 0.64 0.668 ; 
    LAYER M2 ; 
      RECT 3.508 0.576 4.052 0.648 ; 
      RECT 0.076 0.576 2.756 0.648 ; 
      RECT 0.7 0.72 2.108 0.792 ; 
    LAYER V1 ; 
      RECT 3.96 0.576 4.032 0.648 ; 
      RECT 3.528 0.576 3.6 0.648 ; 
      RECT 2.664 0.576 2.736 0.648 ; 
      RECT 2.016 0.72 2.088 0.792 ; 
      RECT 1.584 0.576 1.656 0.648 ; 
      RECT 1.26 0.72 1.332 0.792 ; 
      RECT 0.72 0.72 0.792 0.792 ; 
      RECT 0.568 0.576 0.64 0.648 ; 
      RECT 0.096 0.576 0.168 0.648 ; 
  END 
END DFFHQNx2_ASAP7_75t_R 


MACRO DFFHQNx3_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFHQNx3_ASAP7_75t_R 0 0 ; 
  SIZE 4.752 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.656 0.468 0.944 ; 
        RECT 0.288 0.28 0.468 0.424 ; 
        RECT 0.396 0.136 0.468 0.424 ; 
        RECT 0.288 0.656 0.468 0.8 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.504 1.16 0.576 ; 
        RECT 0.936 0.9 1.084 0.972 ; 
        RECT 0.936 0.108 1.084 0.18 ; 
        RECT 0.936 0.108 1.008 0.972 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.048 0.9 4.684 0.972 ; 
        RECT 4.612 0.108 4.684 0.972 ; 
        RECT 4.048 0.108 4.684 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.752 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.752 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 3.4 0.9 3.816 0.972 ; 
      RECT 3.744 0.108 3.816 0.972 ; 
      RECT 3.096 0.108 3.168 0.476 ; 
      RECT 3.096 0.108 3.816 0.18 ; 
      RECT 2.752 0.896 2.952 0.968 ; 
      RECT 2.88 0.108 2.952 0.968 ; 
      RECT 2.88 0.612 3.6 0.684 ; 
      RECT 3.528 0.468 3.6 0.684 ; 
      RECT 3.312 0.468 3.384 0.684 ; 
      RECT 2.536 0.108 2.952 0.18 ; 
      RECT 2.304 0.9 2.52 0.972 ; 
      RECT 2.448 0.324 2.52 0.972 ; 
      RECT 1.984 0.324 2.52 0.396 ; 
      RECT 2.34 0.18 2.412 0.396 ; 
      RECT 1.456 0.9 1.872 0.972 ; 
      RECT 1.8 0.108 1.872 0.972 ; 
      RECT 1.8 0.488 2.304 0.56 ; 
      RECT 1.672 0.108 1.872 0.18 ; 
      RECT 1.26 0.504 1.332 0.812 ; 
      RECT 1.26 0.504 1.468 0.576 ; 
      RECT 0.592 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.592 0.108 0.792 0.18 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.576 0.188 0.648 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 3.96 0.488 4.032 0.668 ; 
      RECT 2.664 0.404 2.736 0.668 ; 
      RECT 2.016 0.66 2.088 0.812 ; 
      RECT 1.584 0.424 1.656 0.668 ; 
      RECT 0.568 0.424 0.64 0.668 ; 
    LAYER M2 ; 
      RECT 3.508 0.576 4.052 0.648 ; 
      RECT 0.076 0.576 2.756 0.648 ; 
      RECT 0.7 0.72 2.108 0.792 ; 
    LAYER V1 ; 
      RECT 3.96 0.576 4.032 0.648 ; 
      RECT 3.528 0.576 3.6 0.648 ; 
      RECT 2.664 0.576 2.736 0.648 ; 
      RECT 2.016 0.72 2.088 0.792 ; 
      RECT 1.584 0.576 1.656 0.648 ; 
      RECT 1.26 0.72 1.332 0.792 ; 
      RECT 0.72 0.72 0.792 0.792 ; 
      RECT 0.568 0.576 0.64 0.648 ; 
      RECT 0.096 0.576 0.168 0.648 ; 
  END 
END DFFHQNx3_ASAP7_75t_R 


MACRO DFFHQx4_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFHQx4_ASAP7_75t_R 0 0 ; 
  SIZE 5.4 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.656 0.468 0.944 ; 
        RECT 0.288 0.28 0.468 0.424 ; 
        RECT 0.396 0.136 0.468 0.424 ; 
        RECT 0.288 0.656 0.468 0.8 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.504 1.16 0.576 ; 
        RECT 0.936 0.9 1.084 0.972 ; 
        RECT 0.936 0.108 1.084 0.18 ; 
        RECT 0.936 0.108 1.008 0.972 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.5 0.9 5.332 0.972 ; 
        RECT 5.252 0.108 5.332 0.972 ; 
        RECT 4.5 0.108 5.332 0.18 ; 
        RECT 4.5 0.804 4.572 0.972 ; 
        RECT 4.5 0.108 4.572 0.276 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 5.4 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.4 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.048 0.9 4.392 0.972 ; 
      RECT 4.32 0.108 4.392 0.972 ; 
      RECT 4.32 0.508 4.7 0.58 ; 
      RECT 4.048 0.108 4.392 0.18 ; 
      RECT 3.4 0.9 3.816 0.972 ; 
      RECT 3.744 0.108 3.816 0.972 ; 
      RECT 3.096 0.108 3.168 0.476 ; 
      RECT 3.096 0.108 3.816 0.18 ; 
      RECT 2.752 0.896 2.952 0.968 ; 
      RECT 2.88 0.108 2.952 0.968 ; 
      RECT 2.88 0.612 3.6 0.684 ; 
      RECT 3.528 0.468 3.6 0.684 ; 
      RECT 3.312 0.468 3.384 0.684 ; 
      RECT 2.536 0.108 2.952 0.18 ; 
      RECT 2.304 0.9 2.52 0.972 ; 
      RECT 2.448 0.324 2.52 0.972 ; 
      RECT 1.984 0.324 2.52 0.396 ; 
      RECT 2.34 0.18 2.412 0.396 ; 
      RECT 1.456 0.9 1.872 0.972 ; 
      RECT 1.8 0.108 1.872 0.972 ; 
      RECT 1.8 0.488 2.324 0.56 ; 
      RECT 1.672 0.108 1.872 0.18 ; 
      RECT 1.26 0.504 1.332 0.812 ; 
      RECT 1.26 0.504 1.468 0.576 ; 
      RECT 0.592 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.592 0.108 0.792 0.18 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.576 0.188 0.648 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 3.96 0.488 4.032 0.668 ; 
      RECT 2.664 0.404 2.736 0.668 ; 
      RECT 2.016 0.66 2.088 0.812 ; 
      RECT 1.584 0.424 1.656 0.668 ; 
      RECT 0.568 0.424 0.64 0.668 ; 
    LAYER M2 ; 
      RECT 3.508 0.576 4.052 0.648 ; 
      RECT 0.076 0.576 2.756 0.648 ; 
      RECT 0.7 0.72 2.108 0.792 ; 
    LAYER V1 ; 
      RECT 3.96 0.576 4.032 0.648 ; 
      RECT 3.528 0.576 3.6 0.648 ; 
      RECT 2.664 0.576 2.736 0.648 ; 
      RECT 2.016 0.72 2.088 0.792 ; 
      RECT 1.584 0.576 1.656 0.648 ; 
      RECT 1.26 0.72 1.332 0.792 ; 
      RECT 0.72 0.72 0.792 0.792 ; 
      RECT 0.568 0.576 0.64 0.648 ; 
      RECT 0.096 0.576 0.168 0.648 ; 
  END 
END DFFHQx4_ASAP7_75t_R 


MACRO DFFLQNx1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFLQNx1_ASAP7_75t_R 0 0 ; 
  SIZE 4.32 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.656 0.468 0.944 ; 
        RECT 0.288 0.28 0.468 0.424 ; 
        RECT 0.396 0.136 0.468 0.424 ; 
        RECT 0.288 0.656 0.468 0.8 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.9 1.3 0.972 ; 
        RECT 1.152 0.108 1.3 0.18 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.048 0.9 4.248 0.972 ; 
        RECT 4.176 0.108 4.248 0.972 ; 
        RECT 4.048 0.108 4.248 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.32 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.32 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 3.4 0.9 3.816 0.972 ; 
      RECT 3.744 0.108 3.816 0.972 ; 
      RECT 3.096 0.108 3.168 0.476 ; 
      RECT 3.096 0.108 3.816 0.18 ; 
      RECT 2.752 0.9 2.952 0.972 ; 
      RECT 2.88 0.108 2.952 0.972 ; 
      RECT 2.88 0.612 3.6 0.684 ; 
      RECT 3.528 0.468 3.6 0.684 ; 
      RECT 3.312 0.468 3.384 0.684 ; 
      RECT 2.536 0.108 2.952 0.18 ; 
      RECT 2.304 0.9 2.52 0.972 ; 
      RECT 2.448 0.324 2.52 0.972 ; 
      RECT 1.984 0.324 2.52 0.396 ; 
      RECT 2.34 0.136 2.412 0.396 ; 
      RECT 1.456 0.9 1.872 0.972 ; 
      RECT 1.8 0.108 1.872 0.972 ; 
      RECT 1.8 0.488 2.324 0.56 ; 
      RECT 1.672 0.108 1.872 0.18 ; 
      RECT 0.592 0.9 1.008 0.972 ; 
      RECT 0.936 0.108 1.008 0.972 ; 
      RECT 0.592 0.108 1.008 0.18 ; 
      RECT 0.58 0.72 0.792 0.792 ; 
      RECT 0.72 0.504 0.792 0.792 ; 
      RECT 0.484 0.504 0.792 0.576 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.72 0.188 0.792 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 3.96 0.36 4.032 0.668 ; 
      RECT 2.664 0.396 2.736 0.668 ; 
      RECT 2.016 0.66 2.088 0.812 ; 
      RECT 1.584 0.424 1.656 0.668 ; 
      RECT 1.368 0.504 1.44 0.812 ; 
    LAYER M2 ; 
      RECT 3.508 0.576 4.052 0.648 ; 
      RECT 0.916 0.576 2.756 0.648 ; 
      RECT 0.076 0.72 2.108 0.792 ; 
    LAYER V1 ; 
      RECT 3.96 0.576 4.032 0.648 ; 
      RECT 3.528 0.576 3.6 0.648 ; 
      RECT 2.664 0.576 2.736 0.648 ; 
      RECT 2.016 0.72 2.088 0.792 ; 
      RECT 1.584 0.576 1.656 0.648 ; 
      RECT 1.368 0.72 1.44 0.792 ; 
      RECT 0.936 0.576 1.008 0.648 ; 
      RECT 0.6 0.72 0.672 0.792 ; 
      RECT 0.096 0.72 0.168 0.792 ; 
  END 
END DFFLQNx1_ASAP7_75t_R 


MACRO DFFLQNx2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFLQNx2_ASAP7_75t_R 0 0 ; 
  SIZE 4.536 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.048 0.9 4.46 0.972 ; 
        RECT 4.388 0.108 4.46 0.972 ; 
        RECT 4.048 0.108 4.46 0.18 ; 
    END 
  END QN 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.656 0.468 0.944 ; 
        RECT 0.288 0.28 0.468 0.424 ; 
        RECT 0.396 0.136 0.468 0.424 ; 
        RECT 0.288 0.656 0.468 0.8 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.9 1.3 0.972 ; 
        RECT 1.152 0.108 1.3 0.18 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.536 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.536 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 3.4 0.9 3.816 0.972 ; 
      RECT 3.744 0.108 3.816 0.972 ; 
      RECT 3.096 0.108 3.168 0.476 ; 
      RECT 3.096 0.108 3.816 0.18 ; 
      RECT 2.752 0.9 2.952 0.972 ; 
      RECT 2.88 0.108 2.952 0.972 ; 
      RECT 2.88 0.612 3.6 0.684 ; 
      RECT 3.528 0.468 3.6 0.684 ; 
      RECT 3.312 0.468 3.384 0.684 ; 
      RECT 2.536 0.108 2.952 0.18 ; 
      RECT 2.304 0.9 2.52 0.972 ; 
      RECT 2.448 0.324 2.52 0.972 ; 
      RECT 1.984 0.324 2.52 0.396 ; 
      RECT 2.34 0.136 2.412 0.396 ; 
      RECT 1.456 0.9 1.872 0.972 ; 
      RECT 1.8 0.108 1.872 0.972 ; 
      RECT 1.8 0.488 2.324 0.56 ; 
      RECT 1.672 0.108 1.872 0.18 ; 
      RECT 0.592 0.9 1.008 0.972 ; 
      RECT 0.936 0.108 1.008 0.972 ; 
      RECT 0.592 0.108 1.008 0.18 ; 
      RECT 0.58 0.72 0.792 0.792 ; 
      RECT 0.72 0.504 0.792 0.792 ; 
      RECT 0.484 0.504 0.792 0.576 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.72 0.188 0.792 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 3.96 0.36 4.032 0.668 ; 
      RECT 2.664 0.396 2.736 0.668 ; 
      RECT 2.016 0.66 2.088 0.812 ; 
      RECT 1.584 0.424 1.656 0.668 ; 
      RECT 1.368 0.504 1.44 0.812 ; 
    LAYER M2 ; 
      RECT 3.508 0.576 4.052 0.648 ; 
      RECT 0.916 0.576 2.756 0.648 ; 
      RECT 0.076 0.72 2.108 0.792 ; 
    LAYER V1 ; 
      RECT 3.96 0.576 4.032 0.648 ; 
      RECT 3.528 0.576 3.6 0.648 ; 
      RECT 2.664 0.576 2.736 0.648 ; 
      RECT 2.016 0.72 2.088 0.792 ; 
      RECT 1.584 0.576 1.656 0.648 ; 
      RECT 1.368 0.72 1.44 0.792 ; 
      RECT 0.936 0.576 1.008 0.648 ; 
      RECT 0.6 0.72 0.672 0.792 ; 
      RECT 0.096 0.72 0.168 0.792 ; 
  END 
END DFFLQNx2_ASAP7_75t_R 


MACRO DFFLQNx3_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFLQNx3_ASAP7_75t_R 0 0 ; 
  SIZE 4.752 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.656 0.468 0.944 ; 
        RECT 0.288 0.28 0.468 0.424 ; 
        RECT 0.396 0.136 0.468 0.424 ; 
        RECT 0.288 0.656 0.468 0.8 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.9 1.3 0.972 ; 
        RECT 1.152 0.108 1.3 0.18 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.048 0.9 4.684 0.972 ; 
        RECT 4.612 0.108 4.684 0.972 ; 
        RECT 4.044 0.108 4.684 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.752 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.752 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 3.4 0.9 3.816 0.972 ; 
      RECT 3.744 0.108 3.816 0.972 ; 
      RECT 3.096 0.108 3.168 0.476 ; 
      RECT 3.096 0.108 3.816 0.18 ; 
      RECT 2.752 0.9 2.952 0.972 ; 
      RECT 2.88 0.108 2.952 0.972 ; 
      RECT 2.88 0.612 3.6 0.684 ; 
      RECT 3.528 0.468 3.6 0.684 ; 
      RECT 3.312 0.468 3.384 0.684 ; 
      RECT 2.536 0.108 2.952 0.18 ; 
      RECT 2.304 0.9 2.52 0.972 ; 
      RECT 2.448 0.324 2.52 0.972 ; 
      RECT 1.984 0.324 2.52 0.396 ; 
      RECT 2.34 0.136 2.412 0.396 ; 
      RECT 1.456 0.9 1.872 0.972 ; 
      RECT 1.8 0.108 1.872 0.972 ; 
      RECT 1.8 0.488 2.324 0.56 ; 
      RECT 1.672 0.108 1.872 0.18 ; 
      RECT 0.592 0.9 1.008 0.972 ; 
      RECT 0.936 0.108 1.008 0.972 ; 
      RECT 0.592 0.108 1.008 0.18 ; 
      RECT 0.58 0.72 0.792 0.792 ; 
      RECT 0.72 0.504 0.792 0.792 ; 
      RECT 0.484 0.504 0.792 0.576 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.72 0.188 0.792 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 3.96 0.36 4.032 0.668 ; 
      RECT 2.664 0.396 2.736 0.668 ; 
      RECT 2.016 0.66 2.088 0.812 ; 
      RECT 1.584 0.424 1.656 0.668 ; 
      RECT 1.368 0.504 1.44 0.812 ; 
    LAYER M2 ; 
      RECT 3.508 0.576 4.052 0.648 ; 
      RECT 0.916 0.576 2.756 0.648 ; 
      RECT 0.076 0.72 2.108 0.792 ; 
    LAYER V1 ; 
      RECT 3.96 0.576 4.032 0.648 ; 
      RECT 3.528 0.576 3.6 0.648 ; 
      RECT 2.664 0.576 2.736 0.648 ; 
      RECT 2.016 0.72 2.088 0.792 ; 
      RECT 1.584 0.576 1.656 0.648 ; 
      RECT 1.368 0.72 1.44 0.792 ; 
      RECT 0.936 0.576 1.008 0.648 ; 
      RECT 0.6 0.72 0.672 0.792 ; 
      RECT 0.096 0.72 0.168 0.792 ; 
  END 
END DFFLQNx3_ASAP7_75t_R 


MACRO DFFLQx4_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DFFLQx4_ASAP7_75t_R 0 0 ; 
  SIZE 5.4 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.656 0.468 0.944 ; 
        RECT 0.288 0.28 0.468 0.424 ; 
        RECT 0.396 0.136 0.468 0.424 ; 
        RECT 0.288 0.656 0.468 0.8 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.9 1.3 0.972 ; 
        RECT 1.152 0.108 1.3 0.18 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.5 0.9 5.332 0.972 ; 
        RECT 5.252 0.108 5.332 0.972 ; 
        RECT 4.5 0.108 5.332 0.18 ; 
        RECT 4.5 0.804 4.572 0.972 ; 
        RECT 4.5 0.108 4.572 0.276 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 5.4 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.4 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.048 0.9 4.392 0.972 ; 
      RECT 4.32 0.108 4.392 0.972 ; 
      RECT 4.32 0.508 4.7 0.58 ; 
      RECT 4.048 0.108 4.392 0.18 ; 
      RECT 3.4 0.9 3.816 0.972 ; 
      RECT 3.744 0.108 3.816 0.972 ; 
      RECT 3.096 0.108 3.168 0.476 ; 
      RECT 3.096 0.108 3.816 0.18 ; 
      RECT 2.752 0.9 2.952 0.972 ; 
      RECT 2.88 0.108 2.952 0.972 ; 
      RECT 2.88 0.612 3.6 0.684 ; 
      RECT 3.528 0.468 3.6 0.684 ; 
      RECT 3.312 0.468 3.384 0.684 ; 
      RECT 2.536 0.108 2.952 0.18 ; 
      RECT 2.304 0.9 2.52 0.972 ; 
      RECT 2.448 0.324 2.52 0.972 ; 
      RECT 1.984 0.324 2.52 0.396 ; 
      RECT 2.34 0.136 2.412 0.396 ; 
      RECT 1.456 0.9 1.872 0.972 ; 
      RECT 1.8 0.108 1.872 0.972 ; 
      RECT 1.8 0.488 2.324 0.56 ; 
      RECT 1.672 0.108 1.872 0.18 ; 
      RECT 0.592 0.9 1.008 0.972 ; 
      RECT 0.936 0.108 1.008 0.972 ; 
      RECT 0.592 0.108 1.008 0.18 ; 
      RECT 0.58 0.72 0.792 0.792 ; 
      RECT 0.72 0.504 0.792 0.792 ; 
      RECT 0.484 0.504 0.792 0.576 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.72 0.188 0.792 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 3.96 0.488 4.032 0.668 ; 
      RECT 2.664 0.396 2.736 0.668 ; 
      RECT 2.016 0.66 2.088 0.812 ; 
      RECT 1.584 0.424 1.656 0.668 ; 
      RECT 1.368 0.504 1.44 0.812 ; 
    LAYER M2 ; 
      RECT 3.508 0.576 4.052 0.648 ; 
      RECT 0.916 0.576 2.756 0.648 ; 
      RECT 0.076 0.72 2.108 0.792 ; 
    LAYER V1 ; 
      RECT 3.96 0.576 4.032 0.648 ; 
      RECT 3.528 0.576 3.6 0.648 ; 
      RECT 2.664 0.576 2.736 0.648 ; 
      RECT 2.016 0.72 2.088 0.792 ; 
      RECT 1.584 0.576 1.656 0.648 ; 
      RECT 1.368 0.72 1.44 0.792 ; 
      RECT 0.936 0.576 1.008 0.648 ; 
      RECT 0.6 0.72 0.672 0.792 ; 
      RECT 0.096 0.72 0.168 0.792 ; 
  END 
END DFFLQx4_ASAP7_75t_R 


MACRO DHLx1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DHLx1_ASAP7_75t_R 0 0 ; 
  SIZE 3.24 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.612 0.468 0.944 ; 
        RECT 0.288 0.324 0.468 0.468 ; 
        RECT 0.396 0.136 0.468 0.468 ; 
        RECT 0.288 0.612 0.468 0.756 ; 
        RECT 0.288 0.324 0.36 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.108 1.3 0.18 ; 
        RECT 1.152 0.108 1.224 0.944 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.968 0.9 3.168 0.972 ; 
        RECT 3.096 0.108 3.168 0.972 ; 
        RECT 2.968 0.108 3.168 0.18 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.24 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.24 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.32 0.9 2.52 0.972 ; 
      RECT 2.448 0.108 2.52 0.972 ; 
      RECT 2.016 0.108 2.088 0.384 ; 
      RECT 2.016 0.108 2.52 0.18 ; 
      RECT 1.456 0.9 1.872 0.972 ; 
      RECT 1.8 0.108 1.872 0.972 ; 
      RECT 1.8 0.484 2.324 0.556 ; 
      RECT 1.656 0.108 1.872 0.18 ; 
      RECT 1.368 0.756 1.516 0.828 ; 
      RECT 1.368 0.424 1.44 0.828 ; 
      RECT 0.592 0.9 1.008 0.972 ; 
      RECT 0.936 0.108 1.008 0.972 ; 
      RECT 0.592 0.108 1.008 0.18 ; 
      RECT 0.592 0.72 0.792 0.792 ; 
      RECT 0.72 0.504 0.792 0.792 ; 
      RECT 0.552 0.504 0.792 0.576 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.72 0.188 0.792 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 2.88 0.488 2.952 0.668 ; 
      RECT 2.016 0.656 2.088 0.828 ; 
      RECT 1.584 0.424 1.656 0.684 ; 
    LAYER M2 ; 
      RECT 1.8 0.576 2.972 0.648 ; 
      RECT 0.076 0.72 2.108 0.792 ; 
      RECT 0.916 0.576 1.656 0.648 ; 
    LAYER V1 ; 
      RECT 2.88 0.576 2.952 0.648 ; 
      RECT 2.016 0.72 2.088 0.792 ; 
      RECT 1.8 0.576 1.872 0.648 ; 
      RECT 1.584 0.576 1.656 0.648 ; 
      RECT 1.368 0.72 1.44 0.792 ; 
      RECT 0.936 0.576 1.008 0.648 ; 
      RECT 0.612 0.72 0.684 0.792 ; 
      RECT 0.096 0.72 0.168 0.792 ; 
  END 
END DHLx1_ASAP7_75t_R 


MACRO DHLx2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DHLx2_ASAP7_75t_R 0 0 ; 
  SIZE 3.456 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.612 0.468 0.944 ; 
        RECT 0.288 0.324 0.468 0.468 ; 
        RECT 0.396 0.136 0.468 0.468 ; 
        RECT 0.288 0.612 0.468 0.756 ; 
        RECT 0.288 0.324 0.36 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.108 1.3 0.18 ; 
        RECT 1.152 0.108 1.224 0.944 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.964 0.864 3.4 0.936 ; 
        RECT 3.328 0.144 3.4 0.936 ; 
        RECT 2.968 0.144 3.4 0.216 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.456 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.456 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.32 0.9 2.52 0.972 ; 
      RECT 2.448 0.108 2.52 0.972 ; 
      RECT 2.016 0.108 2.088 0.384 ; 
      RECT 2.016 0.108 2.52 0.18 ; 
      RECT 1.456 0.9 1.872 0.972 ; 
      RECT 1.8 0.108 1.872 0.972 ; 
      RECT 1.8 0.484 2.324 0.556 ; 
      RECT 1.656 0.108 1.872 0.18 ; 
      RECT 1.368 0.756 1.516 0.828 ; 
      RECT 1.368 0.424 1.44 0.828 ; 
      RECT 0.592 0.9 1.008 0.972 ; 
      RECT 0.936 0.108 1.008 0.972 ; 
      RECT 0.592 0.108 1.008 0.18 ; 
      RECT 0.592 0.72 0.792 0.792 ; 
      RECT 0.72 0.504 0.792 0.792 ; 
      RECT 0.552 0.504 0.792 0.576 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.72 0.188 0.792 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 3.096 0.36 3.168 0.668 ; 
      RECT 2.88 0.36 2.952 0.668 ; 
      RECT 2.016 0.656 2.088 0.828 ; 
      RECT 1.584 0.424 1.656 0.684 ; 
    LAYER M2 ; 
      RECT 1.8 0.576 3.188 0.648 ; 
      RECT 0.076 0.72 2.108 0.792 ; 
      RECT 0.916 0.576 1.656 0.648 ; 
    LAYER V1 ; 
      RECT 3.096 0.576 3.168 0.648 ; 
      RECT 2.88 0.576 2.952 0.648 ; 
      RECT 2.016 0.72 2.088 0.792 ; 
      RECT 1.8 0.576 1.872 0.648 ; 
      RECT 1.584 0.576 1.656 0.648 ; 
      RECT 1.368 0.72 1.44 0.792 ; 
      RECT 0.936 0.576 1.008 0.648 ; 
      RECT 0.612 0.72 0.684 0.792 ; 
      RECT 0.096 0.72 0.168 0.792 ; 
  END 
END DHLx2_ASAP7_75t_R 


MACRO DHLx3_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DHLx3_ASAP7_75t_R 0 0 ; 
  SIZE 3.672 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.612 0.468 0.944 ; 
        RECT 0.288 0.324 0.468 0.468 ; 
        RECT 0.396 0.136 0.468 0.468 ; 
        RECT 0.288 0.612 0.468 0.756 ; 
        RECT 0.288 0.324 0.36 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.108 1.3 0.18 ; 
        RECT 1.152 0.108 1.224 0.944 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.752 0.9 3.6 0.972 ; 
        RECT 3.528 0.108 3.6 0.972 ; 
        RECT 2.752 0.108 3.6 0.18 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.672 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.672 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.32 0.9 2.52 0.972 ; 
      RECT 2.448 0.108 2.52 0.972 ; 
      RECT 2.016 0.108 2.088 0.384 ; 
      RECT 2.016 0.108 2.52 0.18 ; 
      RECT 1.456 0.9 1.872 0.972 ; 
      RECT 1.8 0.108 1.872 0.972 ; 
      RECT 1.8 0.484 2.324 0.556 ; 
      RECT 1.656 0.108 1.872 0.18 ; 
      RECT 1.368 0.756 1.516 0.828 ; 
      RECT 1.368 0.424 1.44 0.828 ; 
      RECT 0.592 0.9 1.008 0.972 ; 
      RECT 0.936 0.108 1.008 0.972 ; 
      RECT 0.592 0.108 1.008 0.18 ; 
      RECT 0.592 0.72 0.792 0.792 ; 
      RECT 0.72 0.504 0.792 0.792 ; 
      RECT 0.552 0.504 0.792 0.576 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.72 0.188 0.792 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 3.312 0.36 3.384 0.668 ; 
      RECT 3.096 0.36 3.168 0.668 ; 
      RECT 2.88 0.36 2.952 0.668 ; 
      RECT 2.016 0.656 2.088 0.828 ; 
      RECT 1.584 0.424 1.656 0.684 ; 
    LAYER M2 ; 
      RECT 1.8 0.576 3.404 0.648 ; 
      RECT 0.076 0.72 2.108 0.792 ; 
      RECT 0.916 0.576 1.656 0.648 ; 
    LAYER V1 ; 
      RECT 3.312 0.576 3.384 0.648 ; 
      RECT 3.096 0.576 3.168 0.648 ; 
      RECT 2.88 0.576 2.952 0.648 ; 
      RECT 2.016 0.72 2.088 0.792 ; 
      RECT 1.8 0.576 1.872 0.648 ; 
      RECT 1.584 0.576 1.656 0.648 ; 
      RECT 1.368 0.72 1.44 0.792 ; 
      RECT 0.936 0.576 1.008 0.648 ; 
      RECT 0.612 0.72 0.684 0.792 ; 
      RECT 0.096 0.72 0.168 0.792 ; 
  END 
END DHLx3_ASAP7_75t_R 


MACRO DLLx1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DLLx1_ASAP7_75t_R 0 0 ; 
  SIZE 3.24 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.612 0.468 0.944 ; 
        RECT 0.288 0.324 0.468 0.468 ; 
        RECT 0.396 0.136 0.468 0.468 ; 
        RECT 0.288 0.612 0.468 0.756 ; 
        RECT 0.288 0.324 0.36 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.9 1.3 0.972 ; 
        RECT 1.152 0.108 1.3 0.18 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.968 0.9 3.168 0.972 ; 
        RECT 3.096 0.108 3.168 0.972 ; 
        RECT 2.94 0.108 3.168 0.18 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.24 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.24 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.32 0.9 2.52 0.972 ; 
      RECT 2.448 0.108 2.52 0.972 ; 
      RECT 2.016 0.108 2.088 0.388 ; 
      RECT 2.016 0.108 2.52 0.18 ; 
      RECT 1.456 0.9 1.872 0.972 ; 
      RECT 1.8 0.108 1.872 0.972 ; 
      RECT 1.8 0.488 2.32 0.56 ; 
      RECT 1.656 0.108 1.872 0.18 ; 
      RECT 0.592 0.9 1.008 0.972 ; 
      RECT 0.936 0.108 1.008 0.972 ; 
      RECT 0.592 0.108 1.008 0.18 ; 
      RECT 0.592 0.756 0.792 0.828 ; 
      RECT 0.72 0.504 0.792 0.828 ; 
      RECT 0.552 0.504 0.792 0.576 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.576 0.188 0.648 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 2.88 0.424 2.952 0.8 ; 
      RECT 2.016 0.66 2.088 0.812 ; 
      RECT 1.584 0.424 1.656 0.8 ; 
      RECT 1.368 0.424 1.44 0.812 ; 
    LAYER M2 ; 
      RECT 1.8 0.576 2.972 0.648 ; 
      RECT 0.916 0.72 2.108 0.792 ; 
      RECT 0.076 0.576 1.656 0.648 ; 
    LAYER V1 ; 
      RECT 2.88 0.576 2.952 0.648 ; 
      RECT 2.016 0.72 2.088 0.792 ; 
      RECT 1.8 0.576 1.872 0.648 ; 
      RECT 1.584 0.576 1.656 0.648 ; 
      RECT 1.368 0.72 1.44 0.792 ; 
      RECT 0.936 0.72 1.008 0.792 ; 
      RECT 0.72 0.576 0.792 0.648 ; 
      RECT 0.096 0.576 0.168 0.648 ; 
  END 
END DLLx1_ASAP7_75t_R 


MACRO DLLx2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DLLx2_ASAP7_75t_R 0 0 ; 
  SIZE 3.456 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.612 0.468 0.944 ; 
        RECT 0.288 0.324 0.468 0.468 ; 
        RECT 0.396 0.136 0.468 0.468 ; 
        RECT 0.288 0.612 0.468 0.756 ; 
        RECT 0.288 0.324 0.36 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.9 1.3 0.972 ; 
        RECT 1.152 0.108 1.3 0.18 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.752 0.9 3.388 0.972 ; 
        RECT 3.316 0.108 3.388 0.972 ; 
        RECT 2.752 0.108 3.388 0.18 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.456 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.456 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.32 0.9 2.52 0.972 ; 
      RECT 2.448 0.108 2.52 0.972 ; 
      RECT 2.016 0.108 2.088 0.388 ; 
      RECT 2.016 0.108 2.52 0.18 ; 
      RECT 1.456 0.9 1.872 0.972 ; 
      RECT 1.8 0.108 1.872 0.972 ; 
      RECT 1.8 0.488 2.32 0.56 ; 
      RECT 1.656 0.108 1.872 0.18 ; 
      RECT 0.592 0.9 1.008 0.972 ; 
      RECT 0.936 0.108 1.008 0.972 ; 
      RECT 0.592 0.108 1.008 0.18 ; 
      RECT 0.592 0.756 0.792 0.828 ; 
      RECT 0.72 0.504 0.792 0.828 ; 
      RECT 0.552 0.504 0.792 0.576 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.576 0.188 0.648 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 3.096 0.36 3.168 0.668 ; 
      RECT 2.016 0.66 2.088 0.812 ; 
      RECT 1.584 0.424 1.656 0.8 ; 
      RECT 1.368 0.424 1.44 0.812 ; 
    LAYER M2 ; 
      RECT 1.8 0.576 3.2 0.648 ; 
      RECT 0.916 0.72 2.108 0.792 ; 
      RECT 0.076 0.576 1.656 0.648 ; 
    LAYER V1 ; 
      RECT 3.096 0.576 3.168 0.648 ; 
      RECT 2.016 0.72 2.088 0.792 ; 
      RECT 1.8 0.576 1.872 0.648 ; 
      RECT 1.584 0.576 1.656 0.648 ; 
      RECT 1.368 0.72 1.44 0.792 ; 
      RECT 0.936 0.72 1.008 0.792 ; 
      RECT 0.72 0.576 0.792 0.648 ; 
      RECT 0.096 0.576 0.168 0.648 ; 
  END 
END DLLx2_ASAP7_75t_R 


MACRO DLLx3_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN DLLx3_ASAP7_75t_R 0 0 ; 
  SIZE 3.672 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.612 0.468 0.944 ; 
        RECT 0.288 0.324 0.468 0.468 ; 
        RECT 0.396 0.136 0.468 0.468 ; 
        RECT 0.288 0.612 0.468 0.756 ; 
        RECT 0.288 0.324 0.36 0.756 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.9 1.3 0.972 ; 
        RECT 1.152 0.108 1.3 0.18 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
    END 
  END D 
  PIN Q 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.968 0.864 3.604 0.936 ; 
        RECT 3.528 0.144 3.604 0.936 ; 
        RECT 2.968 0.144 3.604 0.216 ; 
    END 
  END Q 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.672 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.672 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 2.32 0.9 2.52 0.972 ; 
      RECT 2.448 0.108 2.52 0.972 ; 
      RECT 2.016 0.108 2.088 0.388 ; 
      RECT 2.016 0.108 2.52 0.18 ; 
      RECT 1.456 0.9 1.872 0.972 ; 
      RECT 1.8 0.108 1.872 0.972 ; 
      RECT 1.8 0.488 2.32 0.56 ; 
      RECT 1.656 0.108 1.872 0.18 ; 
      RECT 0.592 0.9 1.008 0.972 ; 
      RECT 0.936 0.108 1.008 0.972 ; 
      RECT 0.592 0.108 1.008 0.18 ; 
      RECT 0.592 0.756 0.792 0.828 ; 
      RECT 0.72 0.504 0.792 0.828 ; 
      RECT 0.552 0.504 0.792 0.576 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.576 0.188 0.648 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 3.096 0.36 3.168 0.668 ; 
      RECT 2.016 0.66 2.088 0.812 ; 
      RECT 1.584 0.424 1.656 0.8 ; 
      RECT 1.368 0.424 1.44 0.812 ; 
    LAYER M2 ; 
      RECT 1.8 0.576 3.2 0.648 ; 
      RECT 0.916 0.72 2.108 0.792 ; 
      RECT 0.076 0.576 1.656 0.648 ; 
    LAYER V1 ; 
      RECT 3.096 0.576 3.168 0.648 ; 
      RECT 2.016 0.72 2.088 0.792 ; 
      RECT 1.8 0.576 1.872 0.648 ; 
      RECT 1.584 0.576 1.656 0.648 ; 
      RECT 1.368 0.72 1.44 0.792 ; 
      RECT 0.936 0.72 1.008 0.792 ; 
      RECT 0.72 0.576 0.792 0.648 ; 
      RECT 0.096 0.576 0.168 0.648 ; 
  END 
END DLLx3_ASAP7_75t_R 


MACRO FAx1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FAx1_ASAP7_75t_R 0 0 ; 
  SIZE 3.024 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN SN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.296 0.9 1.98 0.972 ; 
        RECT 1.908 0.736 1.98 0.972 ; 
        RECT 1.908 0.108 1.98 0.272 ; 
        RECT 1.296 0.108 1.98 0.18 ; 
        RECT 1.296 0.108 1.368 0.972 ; 
    END 
  END SN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.024 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.236 0.72 2.508 0.792 ; 
      LAYER M1 ; 
        RECT 2.396 0.72 2.52 0.792 ; 
        RECT 2.448 0.484 2.52 0.792 ; 
        RECT 1.532 0.72 1.656 0.792 ; 
        RECT 1.584 0.484 1.656 0.792 ; 
        RECT 0.236 0.72 0.36 0.792 ; 
        RECT 0.288 0.484 0.36 0.792 ; 
      LAYER V1 ; 
        RECT 0.256 0.72 0.328 0.792 ; 
        RECT 1.552 0.72 1.624 0.792 ; 
        RECT 2.416 0.72 2.488 0.792 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.668 0.576 2.756 0.648 ; 
      LAYER M1 ; 
        RECT 2.664 0.484 2.736 0.668 ; 
        RECT 1.152 0.484 1.224 0.668 ; 
        RECT 0.668 0.576 0.792 0.648 ; 
        RECT 0.72 0.484 0.792 0.648 ; 
      LAYER V1 ; 
        RECT 0.688 0.576 0.76 0.648 ; 
        RECT 1.152 0.576 1.224 0.648 ; 
        RECT 2.664 0.576 2.736 0.648 ; 
    END 
  END B 
  PIN CI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.916 0.432 2.348 0.504 ; 
      LAYER M1 ; 
        RECT 2.232 0.432 2.348 0.504 ; 
        RECT 2.232 0.432 2.304 0.596 ; 
        RECT 1.8 0.412 1.872 0.596 ; 
        RECT 0.904 0.432 1.052 0.504 ; 
        RECT 0.936 0.432 1.008 0.596 ; 
      LAYER V1 ; 
        RECT 0.936 0.432 1.008 0.504 ; 
        RECT 1.8 0.432 1.872 0.504 ; 
        RECT 2.256 0.432 2.328 0.504 ; 
    END 
  END CI 
  PIN CON 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.512 0.288 2.172 0.36 ; 
      LAYER M1 ; 
        RECT 2.06 0.288 2.172 0.36 ; 
        RECT 2.016 0.36 2.132 0.432 ; 
        RECT 2.016 0.36 2.088 0.596 ; 
        RECT 0.496 0.288 1.128 0.36 ; 
        RECT 0.496 0.756 0.92 0.828 ; 
        RECT 0.496 0.288 0.568 0.828 ; 
      LAYER V1 ; 
        RECT 0.532 0.288 0.604 0.36 ; 
        RECT 2.08 0.288 2.152 0.36 ; 
    END 
  END CON 
  OBS 
    LAYER M1 ; 
      RECT 2.104 0.108 2.648 0.18 ; 
      RECT 2.104 0.9 2.648 0.972 ; 
      RECT 0.16 0.108 1.136 0.18 ; 
      RECT 0.16 0.9 1.136 0.972 ; 
  END 
END FAx1_ASAP7_75t_R 


MACRO FILLER_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILLER_ASAP7_75t_R 0 0 ; 
  SIZE 0.432 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.432 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.432 0.036 ; 
    END 
  END VSS 
END FILLER_ASAP7_75t_R 


MACRO FILLERxp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN FILLERxp5_ASAP7_75t_R 0 0 ; 
  SIZE 0.216 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.216 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.216 0.036 ; 
    END 
  END VSS 
END FILLERxp5_ASAP7_75t_R 


MACRO HAxp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN HAxp5_ASAP7_75t_R 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.252 1.44 0.6 ; 
        RECT 0.828 0.252 1.44 0.324 ; 
        RECT 0.828 0.108 0.9 0.324 ; 
        RECT 0.072 0.108 0.9 0.18 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.108 0.144 0.944 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.424 0.252 0.576 0.324 ; 
    END 
  END B 
  PIN CON 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.648 0.756 1.656 0.828 ; 
        RECT 1.584 0.484 1.656 0.828 ; 
        RECT 0.376 0.9 0.72 0.972 ; 
        RECT 0.648 0.3 0.72 0.972 ; 
    END 
  END CON 
  PIN SN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.9 1.872 0.972 ; 
        RECT 1.8 0.108 1.872 0.972 ; 
        RECT 1.692 0.108 1.872 0.18 ; 
    END 
  END SN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.944 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 1.024 0.108 1.548 0.18 ; 
  END 
END HAxp5_ASAP7_75t_R 


MACRO HB1xp67_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN HB1xp67_ASAP7_75t_R 0 0 ; 
  SIZE 0.864 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.828 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.864 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.864 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.9 0.792 0.972 ; 
        RECT 0.72 0.108 0.792 0.972 ; 
        RECT 0.592 0.108 0.792 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.468 0.972 ; 
      RECT 0.396 0.612 0.468 0.972 ; 
      RECT 0.396 0.612 0.576 0.684 ; 
      RECT 0.504 0.396 0.576 0.684 ; 
      RECT 0.396 0.396 0.576 0.468 ; 
      RECT 0.396 0.108 0.468 0.468 ; 
      RECT 0.16 0.108 0.468 0.18 ; 
  END 
END HB1xp67_ASAP7_75t_R 


MACRO HB2xp67_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN HB2xp67_ASAP7_75t_R 0 0 ; 
  SIZE 1.08 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.828 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.08 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.9 1.008 0.972 ; 
        RECT 0.936 0.108 1.008 0.972 ; 
        RECT 0.808 0.108 1.008 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.576 0.972 ; 
      RECT 0.504 0.108 0.576 0.972 ; 
      RECT 0.504 0.504 0.812 0.576 ; 
      RECT 0.16 0.108 0.576 0.18 ; 
  END 
END HB2xp67_ASAP7_75t_R 


MACRO HB3xp67_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN HB3xp67_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.828 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.9 1.224 0.972 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
        RECT 1.024 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.72 0.504 1.028 0.576 ; 
      RECT 0.16 0.108 0.792 0.18 ; 
  END 
END HB3xp67_ASAP7_75t_R 


MACRO HB4xp67_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN HB4xp67_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.324 0.22 0.396 ; 
        RECT 0.072 0.324 0.144 0.828 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.24 0.9 1.44 0.972 ; 
        RECT 1.368 0.108 1.44 0.972 ; 
        RECT 1.24 0.108 1.44 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.72 0.504 1.244 0.576 ; 
      RECT 0.16 0.108 0.792 0.18 ; 
  END 
END HB4xp67_ASAP7_75t_R 


MACRO ICGx1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx1_ASAP7_75t_R 0 0 ; 
  SIZE 3.888 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.796 ; 
    END 
  END ENA 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.596 0.9 3.816 0.972 ; 
        RECT 3.744 0.108 3.816 0.972 ; 
        RECT 3.516 0.108 3.816 0.18 ; 
    END 
  END GCLK 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.796 ; 
    END 
  END SE 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.888 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.888 0.036 ; 
    END 
  END VSS 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M2 ; 
        RECT 0.916 0.576 2.54 0.648 ; 
      LAYER M1 ; 
        RECT 2.448 0.712 3.06 0.784 ; 
        RECT 2.988 0.568 3.06 0.784 ; 
        RECT 2.448 0.464 2.52 0.784 ; 
        RECT 1.584 0.576 1.788 0.648 ; 
        RECT 1.584 0.48 1.656 0.648 ; 
        RECT 0.936 0.476 1.008 0.736 ; 
      LAYER V1 ; 
        RECT 0.936 0.576 1.008 0.648 ; 
        RECT 1.656 0.576 1.728 0.648 ; 
        RECT 2.448 0.576 2.52 0.648 ; 
    END 
  END CLK 
  OBS 
    LAYER M1 ; 
      RECT 2.752 0.888 3.384 0.96 ; 
      RECT 3.312 0.752 3.384 0.96 ; 
      RECT 3.312 0.752 3.6 0.824 ; 
      RECT 3.528 0.252 3.6 0.824 ; 
      RECT 2.968 0.252 3.6 0.324 ; 
      RECT 1.024 0.892 1.468 0.964 ; 
      RECT 1.396 0.108 1.468 0.964 ; 
      RECT 1.396 0.724 1.892 0.796 ; 
      RECT 3.312 0.396 3.384 0.588 ; 
      RECT 2.664 0.108 2.736 0.588 ; 
      RECT 2.664 0.396 3.384 0.468 ; 
      RECT 1.24 0.108 2.736 0.18 ; 
      RECT 2.236 0.892 2.436 0.964 ; 
      RECT 2.236 0.308 2.308 0.964 ; 
      RECT 2.236 0.308 2.436 0.38 ; 
      RECT 1.872 0.896 2.088 0.968 ; 
      RECT 2.012 0.292 2.088 0.968 ; 
      RECT 1.568 0.292 2.088 0.364 ; 
      RECT 1.152 0.72 1.296 0.792 ; 
      RECT 1.152 0.288 1.224 0.792 ; 
      RECT 0.148 0.896 0.792 0.968 ; 
      RECT 0.72 0.108 0.792 0.968 ; 
      RECT 0.356 0.108 0.792 0.18 ; 
    LAYER M2 ; 
      RECT 1.184 0.72 2.328 0.792 ; 
    LAYER V1 ; 
      RECT 2.236 0.72 2.308 0.792 ; 
      RECT 1.204 0.72 1.276 0.792 ; 
  END 
END ICGx1_ASAP7_75t_R 


MACRO ICGx2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx2_ASAP7_75t_R 0 0 ; 
  SIZE 4.104 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.796 ; 
    END 
  END ENA 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.596 0.9 4.032 0.972 ; 
        RECT 3.96 0.108 4.032 0.972 ; 
        RECT 3.516 0.108 4.032 0.18 ; 
    END 
  END GCLK 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.796 ; 
    END 
  END SE 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.104 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.104 0.036 ; 
    END 
  END VSS 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M2 ; 
        RECT 0.916 0.576 2.54 0.648 ; 
      LAYER M1 ; 
        RECT 2.448 0.712 3.06 0.784 ; 
        RECT 2.988 0.568 3.06 0.784 ; 
        RECT 2.448 0.464 2.52 0.784 ; 
        RECT 1.584 0.576 1.788 0.648 ; 
        RECT 1.584 0.48 1.656 0.648 ; 
        RECT 0.936 0.476 1.008 0.736 ; 
      LAYER V1 ; 
        RECT 0.936 0.576 1.008 0.648 ; 
        RECT 1.656 0.576 1.728 0.648 ; 
        RECT 2.448 0.576 2.52 0.648 ; 
    END 
  END CLK 
  OBS 
    LAYER M1 ; 
      RECT 2.752 0.888 3.384 0.96 ; 
      RECT 3.312 0.752 3.384 0.96 ; 
      RECT 3.312 0.752 3.6 0.824 ; 
      RECT 3.528 0.252 3.6 0.824 ; 
      RECT 2.968 0.252 3.6 0.324 ; 
      RECT 1.024 0.892 1.468 0.964 ; 
      RECT 1.396 0.108 1.468 0.964 ; 
      RECT 1.396 0.724 1.892 0.796 ; 
      RECT 3.312 0.396 3.384 0.588 ; 
      RECT 2.664 0.108 2.736 0.588 ; 
      RECT 2.664 0.396 3.384 0.468 ; 
      RECT 1.24 0.108 2.736 0.18 ; 
      RECT 2.236 0.892 2.436 0.964 ; 
      RECT 2.236 0.308 2.308 0.964 ; 
      RECT 2.236 0.308 2.436 0.38 ; 
      RECT 1.872 0.896 2.088 0.968 ; 
      RECT 2.012 0.292 2.088 0.968 ; 
      RECT 1.568 0.292 2.088 0.364 ; 
      RECT 1.152 0.72 1.296 0.792 ; 
      RECT 1.152 0.288 1.224 0.792 ; 
      RECT 1.028 0.288 1.224 0.36 ; 
      RECT 0.148 0.896 0.792 0.968 ; 
      RECT 0.72 0.108 0.792 0.968 ; 
      RECT 0.356 0.108 0.792 0.18 ; 
    LAYER M2 ; 
      RECT 1.184 0.72 2.328 0.792 ; 
    LAYER V1 ; 
      RECT 2.236 0.72 2.308 0.792 ; 
      RECT 1.204 0.72 1.276 0.792 ; 
  END 
END ICGx2_ASAP7_75t_R 


MACRO ICGx2p67DC_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx2p67DC_ASAP7_75t_R 0 0 ; 
  SIZE 10.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 9.864 0.9 10.084 0.972 ; 
        RECT 10.012 0.108 10.084 0.972 ; 
        RECT 9.784 0.108 10.084 0.18 ; 
        RECT 7.704 0.9 7.924 0.972 ; 
        RECT 7.852 0.108 7.924 0.972 ; 
        RECT 7.624 0.108 7.924 0.18 ; 
        RECT 2.452 0.108 2.752 0.18 ; 
        RECT 2.452 0.9 2.672 0.972 ; 
        RECT 2.452 0.108 2.524 0.972 ; 
        RECT 0.292 0.108 0.592 0.18 ; 
        RECT 0.292 0.9 0.512 0.972 ; 
        RECT 0.292 0.108 0.364 0.972 ; 
      LAYER M2 ; 
        RECT 0.248 0.144 10.128 0.216 ; 
      LAYER V1 ; 
        RECT 0.292 0.144 0.364 0.216 ; 
        RECT 2.452 0.144 2.524 0.216 ; 
        RECT 7.852 0.144 7.924 0.216 ; 
        RECT 10.012 0.144 10.084 0.216 ; 
    END 
  END GCLK 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 10.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 10.376 0.036 ; 
    END 
  END VSS 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 9.128 0.684 9.404 0.756 ; 
        RECT 9.332 0.54 9.404 0.756 ; 
        RECT 9.172 0.54 9.404 0.612 ; 
        RECT 6.556 0.712 7.168 0.784 ; 
        RECT 7.096 0.568 7.168 0.784 ; 
        RECT 6.556 0.464 6.628 0.784 ; 
        RECT 5.692 0.576 5.896 0.648 ; 
        RECT 5.692 0.48 5.764 0.648 ; 
        RECT 5.044 0.476 5.116 0.736 ; 
        RECT 3.208 0.712 3.82 0.784 ; 
        RECT 3.748 0.464 3.82 0.784 ; 
        RECT 3.208 0.568 3.28 0.784 ; 
        RECT 0.996 0.684 1.272 0.756 ; 
        RECT 0.996 0.54 1.228 0.612 ; 
        RECT 0.996 0.54 1.068 0.756 ; 
      LAYER M2 ; 
        RECT 0.944 0.576 9.436 0.648 ; 
      LAYER V1 ; 
        RECT 0.996 0.576 1.068 0.648 ; 
        RECT 3.748 0.576 3.82 0.648 ; 
        RECT 5.044 0.576 5.116 0.648 ; 
        RECT 5.764 0.576 5.836 0.648 ; 
        RECT 6.556 0.576 6.628 0.648 ; 
        RECT 9.332 0.576 9.404 0.648 ; 
    END 
  END CLK 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.308 0.688 4.468 0.796 ; 
        RECT 4.396 0.28 4.468 0.796 ; 
        RECT 4.132 0.888 4.384 0.964 ; 
        RECT 4.308 0.688 4.384 0.964 ; 
      LAYER M2 ; 
        RECT 3.932 0.864 4.952 0.936 ; 
      LAYER V1 ; 
        RECT 4.308 0.864 4.384 0.936 ; 
    END 
  END ENA 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.612 0.28 4.684 0.796 ; 
      LAYER M2 ; 
        RECT 3.932 0.288 4.952 0.36 ; 
      LAYER V1 ; 
        RECT 4.612 0.288 4.684 0.36 ; 
    END 
  END SE 
  OBS 
    LAYER M1 ; 
      RECT 9.02 0.888 9.652 0.96 ; 
      RECT 9.58 0.752 9.652 0.96 ; 
      RECT 9.58 0.752 9.868 0.824 ; 
      RECT 9.796 0.252 9.868 0.824 ; 
      RECT 9.236 0.252 9.868 0.324 ; 
      RECT 9.58 0.396 9.652 0.588 ; 
      RECT 8.932 0.396 9.004 0.588 ; 
      RECT 8.932 0.396 9.652 0.468 ; 
      RECT 8.5 0.504 8.724 0.576 ; 
      RECT 8.5 0.36 8.572 0.576 ; 
      RECT 8.156 0.36 8.764 0.432 ; 
      RECT 8.08 0.648 8.7 0.72 ; 
      RECT 8.284 0.504 8.356 0.72 ; 
      RECT 8.124 0.504 8.356 0.576 ; 
      RECT 6.86 0.888 7.492 0.96 ; 
      RECT 7.42 0.752 7.492 0.96 ; 
      RECT 7.42 0.752 7.708 0.824 ; 
      RECT 7.636 0.252 7.708 0.824 ; 
      RECT 7.076 0.252 7.708 0.324 ; 
      RECT 5.132 0.892 5.576 0.964 ; 
      RECT 5.504 0.108 5.576 0.964 ; 
      RECT 5.504 0.724 6 0.796 ; 
      RECT 7.42 0.396 7.492 0.588 ; 
      RECT 6.772 0.108 6.844 0.588 ; 
      RECT 6.772 0.396 7.492 0.468 ; 
      RECT 5.348 0.108 6.844 0.18 ; 
      RECT 6.344 0.892 6.544 0.964 ; 
      RECT 6.344 0.308 6.416 0.964 ; 
      RECT 6.344 0.308 6.544 0.38 ; 
      RECT 5.98 0.896 6.196 0.968 ; 
      RECT 6.12 0.292 6.196 0.968 ; 
      RECT 5.676 0.292 6.196 0.364 ; 
      RECT 5.26 0.72 5.404 0.792 ; 
      RECT 5.26 0.288 5.332 0.792 ; 
      RECT 5.136 0.288 5.332 0.36 ; 
      RECT 4.484 0.896 4.9 0.968 ; 
      RECT 4.828 0.108 4.9 0.968 ; 
      RECT 4.464 0.108 4.9 0.18 ; 
      RECT 3.832 0.892 4.032 0.964 ; 
      RECT 3.96 0.308 4.032 0.964 ; 
      RECT 3.832 0.308 4.032 0.38 ; 
      RECT 3.532 0.396 3.604 0.588 ; 
      RECT 2.884 0.396 2.956 0.588 ; 
      RECT 2.884 0.396 3.604 0.468 ; 
      RECT 2.884 0.888 3.516 0.96 ; 
      RECT 2.884 0.752 2.956 0.96 ; 
      RECT 2.668 0.752 2.956 0.824 ; 
      RECT 2.668 0.252 2.74 0.824 ; 
      RECT 2.668 0.252 3.3 0.324 ; 
      RECT 1.676 0.648 2.296 0.72 ; 
      RECT 2.02 0.504 2.092 0.72 ; 
      RECT 2.02 0.504 2.252 0.576 ; 
      RECT 1.652 0.504 1.876 0.576 ; 
      RECT 1.804 0.36 1.876 0.576 ; 
      RECT 1.612 0.36 2.22 0.432 ; 
      RECT 1.372 0.396 1.444 0.588 ; 
      RECT 0.724 0.396 0.796 0.588 ; 
      RECT 0.724 0.396 1.444 0.468 ; 
      RECT 0.724 0.888 1.356 0.96 ; 
      RECT 0.724 0.752 0.796 0.96 ; 
      RECT 0.508 0.752 0.796 0.824 ; 
      RECT 0.508 0.252 0.58 0.824 ; 
      RECT 0.508 0.252 1.14 0.324 ; 
    LAYER M2 ; 
      RECT 1.348 0.432 9.028 0.504 ; 
      RECT 3.932 0.72 6.436 0.792 ; 
    LAYER V1 ; 
      RECT 8.932 0.432 9.004 0.504 ; 
      RECT 6.772 0.432 6.844 0.504 ; 
      RECT 6.344 0.72 6.416 0.792 ; 
      RECT 5.312 0.72 5.384 0.792 ; 
      RECT 3.96 0.72 4.032 0.792 ; 
      RECT 3.532 0.432 3.604 0.504 ; 
      RECT 1.372 0.432 1.444 0.504 ; 
  END 
END ICGx2p67DC_ASAP7_75t_R 


MACRO ICGx3_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx3_ASAP7_75t_R 0 0 ; 
  SIZE 4.32 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.796 ; 
    END 
  END ENA 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.596 0.9 4.248 0.972 ; 
        RECT 4.176 0.108 4.248 0.972 ; 
        RECT 3.516 0.108 4.248 0.18 ; 
    END 
  END GCLK 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.796 ; 
    END 
  END SE 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.32 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.32 0.036 ; 
    END 
  END VSS 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M2 ; 
        RECT 0.916 0.576 2.54 0.648 ; 
      LAYER M1 ; 
        RECT 2.448 0.712 3.06 0.784 ; 
        RECT 2.988 0.568 3.06 0.784 ; 
        RECT 2.448 0.464 2.52 0.784 ; 
        RECT 1.584 0.576 1.788 0.648 ; 
        RECT 1.584 0.48 1.656 0.648 ; 
        RECT 0.936 0.476 1.008 0.736 ; 
      LAYER V1 ; 
        RECT 0.936 0.576 1.008 0.648 ; 
        RECT 1.656 0.576 1.728 0.648 ; 
        RECT 2.448 0.576 2.52 0.648 ; 
    END 
  END CLK 
  OBS 
    LAYER M1 ; 
      RECT 2.752 0.888 3.384 0.96 ; 
      RECT 3.312 0.752 3.384 0.96 ; 
      RECT 3.312 0.752 3.6 0.824 ; 
      RECT 3.528 0.252 3.6 0.824 ; 
      RECT 2.968 0.252 3.6 0.324 ; 
      RECT 1.024 0.892 1.468 0.964 ; 
      RECT 1.396 0.108 1.468 0.964 ; 
      RECT 1.396 0.724 1.892 0.796 ; 
      RECT 3.312 0.396 3.384 0.588 ; 
      RECT 2.664 0.108 2.736 0.588 ; 
      RECT 2.664 0.396 3.384 0.468 ; 
      RECT 1.24 0.108 2.736 0.18 ; 
      RECT 2.236 0.892 2.436 0.964 ; 
      RECT 2.236 0.308 2.308 0.964 ; 
      RECT 2.236 0.308 2.436 0.38 ; 
      RECT 1.872 0.896 2.088 0.968 ; 
      RECT 2.012 0.292 2.088 0.968 ; 
      RECT 1.568 0.292 2.088 0.364 ; 
      RECT 1.152 0.72 1.296 0.792 ; 
      RECT 1.152 0.288 1.224 0.792 ; 
      RECT 1.028 0.288 1.224 0.36 ; 
      RECT 0.148 0.896 0.792 0.968 ; 
      RECT 0.72 0.108 0.792 0.968 ; 
      RECT 0.356 0.108 0.792 0.18 ; 
    LAYER M2 ; 
      RECT 1.184 0.72 2.328 0.792 ; 
    LAYER V1 ; 
      RECT 2.236 0.72 2.308 0.792 ; 
      RECT 1.204 0.72 1.276 0.792 ; 
  END 
END ICGx3_ASAP7_75t_R 


MACRO ICGx4DC_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx4DC_ASAP7_75t_R 0 0 ; 
  SIZE 10.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 9.864 0.9 10.084 0.972 ; 
        RECT 10.012 0.108 10.084 0.972 ; 
        RECT 9.784 0.108 10.084 0.18 ; 
        RECT 7.704 0.9 7.924 0.972 ; 
        RECT 7.852 0.108 7.924 0.972 ; 
        RECT 7.624 0.108 7.924 0.18 ; 
        RECT 2.452 0.108 2.752 0.18 ; 
        RECT 2.452 0.9 2.672 0.972 ; 
        RECT 2.452 0.108 2.524 0.972 ; 
        RECT 0.292 0.108 0.592 0.18 ; 
        RECT 0.292 0.9 0.512 0.972 ; 
        RECT 0.292 0.108 0.364 0.972 ; 
      LAYER M2 ; 
        RECT 0.248 0.144 10.128 0.216 ; 
      LAYER V1 ; 
        RECT 0.292 0.144 0.364 0.216 ; 
        RECT 2.452 0.144 2.524 0.216 ; 
        RECT 7.852 0.144 7.924 0.216 ; 
        RECT 10.012 0.144 10.084 0.216 ; 
    END 
  END GCLK 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 10.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 10.376 0.036 ; 
    END 
  END VSS 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 9.128 0.684 9.404 0.756 ; 
        RECT 9.332 0.54 9.404 0.756 ; 
        RECT 9.172 0.54 9.404 0.612 ; 
        RECT 6.556 0.712 7.168 0.784 ; 
        RECT 7.096 0.568 7.168 0.784 ; 
        RECT 6.556 0.464 6.628 0.784 ; 
        RECT 5.692 0.576 5.896 0.648 ; 
        RECT 5.692 0.48 5.764 0.648 ; 
        RECT 5.044 0.476 5.116 0.736 ; 
        RECT 3.208 0.712 3.82 0.784 ; 
        RECT 3.748 0.464 3.82 0.784 ; 
        RECT 3.208 0.568 3.28 0.784 ; 
        RECT 0.996 0.684 1.272 0.756 ; 
        RECT 0.996 0.54 1.228 0.612 ; 
        RECT 0.996 0.54 1.068 0.756 ; 
      LAYER M2 ; 
        RECT 0.944 0.576 9.436 0.648 ; 
      LAYER V1 ; 
        RECT 0.996 0.576 1.068 0.648 ; 
        RECT 3.748 0.576 3.82 0.648 ; 
        RECT 5.044 0.576 5.116 0.648 ; 
        RECT 5.764 0.576 5.836 0.648 ; 
        RECT 6.556 0.576 6.628 0.648 ; 
        RECT 9.332 0.576 9.404 0.648 ; 
    END 
  END CLK 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.308 0.688 4.468 0.796 ; 
        RECT 4.396 0.28 4.468 0.796 ; 
        RECT 4.132 0.888 4.384 0.964 ; 
        RECT 4.308 0.688 4.384 0.964 ; 
      LAYER M2 ; 
        RECT 3.932 0.864 4.952 0.936 ; 
      LAYER V1 ; 
        RECT 4.308 0.864 4.384 0.936 ; 
    END 
  END ENA 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.612 0.28 4.684 0.796 ; 
      LAYER M2 ; 
        RECT 3.932 0.288 4.952 0.36 ; 
      LAYER V1 ; 
        RECT 4.612 0.288 4.684 0.36 ; 
    END 
  END SE 
  OBS 
    LAYER M1 ; 
      RECT 9.02 0.888 9.652 0.96 ; 
      RECT 9.58 0.752 9.652 0.96 ; 
      RECT 9.58 0.752 9.868 0.824 ; 
      RECT 9.796 0.252 9.868 0.824 ; 
      RECT 9.236 0.252 9.868 0.324 ; 
      RECT 9.58 0.396 9.652 0.588 ; 
      RECT 8.932 0.396 9.004 0.588 ; 
      RECT 8.932 0.396 9.652 0.468 ; 
      RECT 8.5 0.504 8.724 0.576 ; 
      RECT 8.5 0.36 8.572 0.576 ; 
      RECT 8.156 0.36 8.764 0.432 ; 
      RECT 8.08 0.648 8.7 0.72 ; 
      RECT 8.284 0.504 8.356 0.72 ; 
      RECT 8.124 0.504 8.356 0.576 ; 
      RECT 6.86 0.888 7.492 0.96 ; 
      RECT 7.42 0.752 7.492 0.96 ; 
      RECT 7.42 0.752 7.708 0.824 ; 
      RECT 7.636 0.252 7.708 0.824 ; 
      RECT 7.076 0.252 7.708 0.324 ; 
      RECT 5.132 0.892 5.576 0.964 ; 
      RECT 5.504 0.108 5.576 0.964 ; 
      RECT 5.504 0.724 6 0.796 ; 
      RECT 7.42 0.396 7.492 0.588 ; 
      RECT 6.772 0.108 6.844 0.588 ; 
      RECT 6.772 0.396 7.492 0.468 ; 
      RECT 5.348 0.108 6.844 0.18 ; 
      RECT 6.344 0.892 6.544 0.964 ; 
      RECT 6.344 0.308 6.416 0.964 ; 
      RECT 6.344 0.308 6.544 0.38 ; 
      RECT 5.98 0.896 6.196 0.968 ; 
      RECT 6.12 0.292 6.196 0.968 ; 
      RECT 5.676 0.292 6.196 0.364 ; 
      RECT 5.26 0.72 5.404 0.792 ; 
      RECT 5.26 0.288 5.332 0.792 ; 
      RECT 5.136 0.288 5.332 0.36 ; 
      RECT 4.484 0.896 4.9 0.968 ; 
      RECT 4.828 0.108 4.9 0.968 ; 
      RECT 4.464 0.108 4.9 0.18 ; 
      RECT 3.832 0.892 4.032 0.964 ; 
      RECT 3.96 0.308 4.032 0.964 ; 
      RECT 3.832 0.308 4.032 0.38 ; 
      RECT 3.532 0.396 3.604 0.588 ; 
      RECT 2.884 0.396 2.956 0.588 ; 
      RECT 2.884 0.396 3.604 0.468 ; 
      RECT 2.884 0.888 3.516 0.96 ; 
      RECT 2.884 0.752 2.956 0.96 ; 
      RECT 2.668 0.752 2.956 0.824 ; 
      RECT 2.668 0.252 2.74 0.824 ; 
      RECT 2.668 0.252 3.3 0.324 ; 
      RECT 1.676 0.648 2.296 0.72 ; 
      RECT 2.02 0.504 2.092 0.72 ; 
      RECT 2.02 0.504 2.252 0.576 ; 
      RECT 1.652 0.504 1.876 0.576 ; 
      RECT 1.804 0.36 1.876 0.576 ; 
      RECT 1.612 0.36 2.22 0.432 ; 
      RECT 1.372 0.396 1.444 0.588 ; 
      RECT 0.724 0.396 0.796 0.588 ; 
      RECT 0.724 0.396 1.444 0.468 ; 
      RECT 0.724 0.888 1.356 0.96 ; 
      RECT 0.724 0.752 0.796 0.96 ; 
      RECT 0.508 0.752 0.796 0.824 ; 
      RECT 0.508 0.252 0.58 0.824 ; 
      RECT 0.508 0.252 1.14 0.324 ; 
    LAYER M2 ; 
      RECT 1.348 0.432 9.028 0.504 ; 
      RECT 3.932 0.72 6.436 0.792 ; 
    LAYER V1 ; 
      RECT 8.932 0.432 9.004 0.504 ; 
      RECT 6.772 0.432 6.844 0.504 ; 
      RECT 6.344 0.72 6.416 0.792 ; 
      RECT 5.312 0.72 5.384 0.792 ; 
      RECT 3.96 0.72 4.032 0.792 ; 
      RECT 3.532 0.432 3.604 0.504 ; 
      RECT 1.372 0.432 1.444 0.504 ; 
  END 
END ICGx4DC_ASAP7_75t_R 


MACRO ICGx4_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx4_ASAP7_75t_R 0 0 ; 
  SIZE 4.536 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.796 ; 
    END 
  END ENA 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.56 0.9 4.248 0.972 ; 
        RECT 4.176 0.108 4.248 0.972 ; 
        RECT 3.556 0.108 4.248 0.18 ; 
    END 
  END GCLK 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.796 ; 
    END 
  END SE 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.536 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.536 0.036 ; 
    END 
  END VSS 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M2 ; 
        RECT 0.916 0.576 2.54 0.648 ; 
      LAYER M1 ; 
        RECT 2.448 0.712 3.06 0.784 ; 
        RECT 2.988 0.568 3.06 0.784 ; 
        RECT 2.448 0.464 2.52 0.784 ; 
        RECT 1.584 0.576 1.788 0.648 ; 
        RECT 1.584 0.48 1.656 0.648 ; 
        RECT 0.936 0.476 1.008 0.736 ; 
      LAYER V1 ; 
        RECT 0.936 0.576 1.008 0.648 ; 
        RECT 1.656 0.576 1.728 0.648 ; 
        RECT 2.448 0.576 2.52 0.648 ; 
    END 
  END CLK 
  OBS 
    LAYER M1 ; 
      RECT 2.752 0.888 3.384 0.96 ; 
      RECT 3.312 0.752 3.384 0.96 ; 
      RECT 3.312 0.752 3.6 0.824 ; 
      RECT 3.528 0.252 3.6 0.824 ; 
      RECT 2.968 0.252 3.6 0.324 ; 
      RECT 1.024 0.892 1.468 0.964 ; 
      RECT 1.396 0.108 1.468 0.964 ; 
      RECT 1.396 0.724 1.892 0.796 ; 
      RECT 3.312 0.396 3.384 0.588 ; 
      RECT 2.664 0.108 2.736 0.588 ; 
      RECT 2.664 0.396 3.384 0.468 ; 
      RECT 1.24 0.108 2.736 0.18 ; 
      RECT 2.236 0.892 2.436 0.964 ; 
      RECT 2.236 0.308 2.308 0.964 ; 
      RECT 2.236 0.308 2.436 0.38 ; 
      RECT 1.872 0.896 2.088 0.968 ; 
      RECT 2.012 0.292 2.088 0.968 ; 
      RECT 1.568 0.292 2.088 0.364 ; 
      RECT 1.152 0.72 1.296 0.792 ; 
      RECT 1.152 0.288 1.224 0.792 ; 
      RECT 1.028 0.288 1.224 0.36 ; 
      RECT 0.148 0.896 0.792 0.968 ; 
      RECT 0.72 0.108 0.792 0.968 ; 
      RECT 0.356 0.108 0.792 0.18 ; 
    LAYER M2 ; 
      RECT 1.184 0.72 2.328 0.792 ; 
    LAYER V1 ; 
      RECT 2.236 0.72 2.308 0.792 ; 
      RECT 1.204 0.72 1.276 0.792 ; 
  END 
END ICGx4_ASAP7_75t_R 


MACRO ICGx5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx5_ASAP7_75t_R 0 0 ; 
  SIZE 4.752 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.796 ; 
    END 
  END ENA 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.56 0.9 4.68 0.972 ; 
        RECT 4.608 0.108 4.68 0.972 ; 
        RECT 3.556 0.108 4.68 0.18 ; 
    END 
  END GCLK 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.796 ; 
    END 
  END SE 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.752 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.752 0.036 ; 
    END 
  END VSS 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M2 ; 
        RECT 0.916 0.576 2.54 0.648 ; 
      LAYER M1 ; 
        RECT 2.448 0.712 3.06 0.784 ; 
        RECT 2.988 0.568 3.06 0.784 ; 
        RECT 2.448 0.464 2.52 0.784 ; 
        RECT 1.584 0.576 1.788 0.648 ; 
        RECT 1.584 0.48 1.656 0.648 ; 
        RECT 0.936 0.476 1.008 0.736 ; 
      LAYER V1 ; 
        RECT 0.936 0.576 1.008 0.648 ; 
        RECT 1.656 0.576 1.728 0.648 ; 
        RECT 2.448 0.576 2.52 0.648 ; 
    END 
  END CLK 
  OBS 
    LAYER M1 ; 
      RECT 2.752 0.888 3.384 0.96 ; 
      RECT 3.312 0.752 3.384 0.96 ; 
      RECT 3.312 0.752 3.6 0.824 ; 
      RECT 3.528 0.252 3.6 0.824 ; 
      RECT 2.968 0.252 3.6 0.324 ; 
      RECT 1.024 0.892 1.468 0.964 ; 
      RECT 1.396 0.108 1.468 0.964 ; 
      RECT 1.396 0.724 1.892 0.796 ; 
      RECT 3.312 0.396 3.384 0.588 ; 
      RECT 2.664 0.108 2.736 0.588 ; 
      RECT 2.664 0.396 3.384 0.468 ; 
      RECT 1.24 0.108 2.736 0.18 ; 
      RECT 2.236 0.892 2.436 0.964 ; 
      RECT 2.236 0.308 2.308 0.964 ; 
      RECT 2.236 0.308 2.436 0.38 ; 
      RECT 1.872 0.896 2.088 0.968 ; 
      RECT 2.012 0.292 2.088 0.968 ; 
      RECT 1.568 0.292 2.088 0.364 ; 
      RECT 1.152 0.72 1.296 0.792 ; 
      RECT 1.152 0.288 1.224 0.792 ; 
      RECT 1.028 0.288 1.224 0.36 ; 
      RECT 0.148 0.896 0.792 0.968 ; 
      RECT 0.72 0.108 0.792 0.968 ; 
      RECT 0.356 0.108 0.792 0.18 ; 
    LAYER M2 ; 
      RECT 1.184 0.72 2.328 0.792 ; 
    LAYER V1 ; 
      RECT 2.236 0.72 2.308 0.792 ; 
      RECT 1.204 0.72 1.276 0.792 ; 
  END 
END ICGx5_ASAP7_75t_R 


MACRO ICGx5p33DC_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx5p33DC_ASAP7_75t_R 0 0 ; 
  SIZE 10.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 9.864 0.9 10.084 0.972 ; 
        RECT 10.012 0.108 10.084 0.972 ; 
        RECT 9.784 0.108 10.084 0.18 ; 
        RECT 7.704 0.9 7.924 0.972 ; 
        RECT 7.852 0.108 7.924 0.972 ; 
        RECT 7.624 0.108 7.924 0.18 ; 
        RECT 2.452 0.108 2.752 0.18 ; 
        RECT 2.452 0.9 2.672 0.972 ; 
        RECT 2.452 0.108 2.524 0.972 ; 
        RECT 0.292 0.108 0.592 0.18 ; 
        RECT 0.292 0.9 0.512 0.972 ; 
        RECT 0.292 0.108 0.364 0.972 ; 
      LAYER M2 ; 
        RECT 0.248 0.144 10.128 0.216 ; 
      LAYER V1 ; 
        RECT 0.292 0.144 0.364 0.216 ; 
        RECT 2.452 0.144 2.524 0.216 ; 
        RECT 7.852 0.144 7.924 0.216 ; 
        RECT 10.012 0.144 10.084 0.216 ; 
    END 
  END GCLK 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 10.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 10.376 0.036 ; 
    END 
  END VSS 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 9.128 0.684 9.404 0.756 ; 
        RECT 9.332 0.54 9.404 0.756 ; 
        RECT 9.172 0.54 9.404 0.612 ; 
        RECT 6.556 0.712 7.168 0.784 ; 
        RECT 7.096 0.568 7.168 0.784 ; 
        RECT 6.556 0.464 6.628 0.784 ; 
        RECT 5.692 0.576 5.896 0.648 ; 
        RECT 5.692 0.48 5.764 0.648 ; 
        RECT 5.044 0.476 5.116 0.736 ; 
        RECT 3.208 0.712 3.82 0.784 ; 
        RECT 3.748 0.464 3.82 0.784 ; 
        RECT 3.208 0.568 3.28 0.784 ; 
        RECT 0.996 0.684 1.272 0.756 ; 
        RECT 0.996 0.54 1.228 0.612 ; 
        RECT 0.996 0.54 1.068 0.756 ; 
      LAYER M2 ; 
        RECT 0.944 0.576 9.436 0.648 ; 
      LAYER V1 ; 
        RECT 0.996 0.576 1.068 0.648 ; 
        RECT 3.748 0.576 3.82 0.648 ; 
        RECT 5.044 0.576 5.116 0.648 ; 
        RECT 5.764 0.576 5.836 0.648 ; 
        RECT 6.556 0.576 6.628 0.648 ; 
        RECT 9.332 0.576 9.404 0.648 ; 
    END 
  END CLK 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.308 0.688 4.468 0.796 ; 
        RECT 4.396 0.28 4.468 0.796 ; 
        RECT 4.132 0.888 4.384 0.964 ; 
        RECT 4.308 0.688 4.384 0.964 ; 
      LAYER M2 ; 
        RECT 3.932 0.864 4.952 0.936 ; 
      LAYER V1 ; 
        RECT 4.308 0.864 4.384 0.936 ; 
    END 
  END ENA 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.612 0.28 4.684 0.796 ; 
      LAYER M2 ; 
        RECT 3.932 0.288 4.952 0.36 ; 
      LAYER V1 ; 
        RECT 4.612 0.288 4.684 0.36 ; 
    END 
  END SE 
  OBS 
    LAYER M1 ; 
      RECT 9.02 0.888 9.652 0.96 ; 
      RECT 9.58 0.752 9.652 0.96 ; 
      RECT 9.58 0.752 9.868 0.824 ; 
      RECT 9.796 0.252 9.868 0.824 ; 
      RECT 9.236 0.252 9.868 0.324 ; 
      RECT 9.58 0.396 9.652 0.588 ; 
      RECT 8.932 0.396 9.004 0.588 ; 
      RECT 8.932 0.396 9.652 0.468 ; 
      RECT 8.5 0.504 8.724 0.576 ; 
      RECT 8.5 0.36 8.572 0.576 ; 
      RECT 8.156 0.36 8.764 0.432 ; 
      RECT 8.08 0.648 8.7 0.72 ; 
      RECT 8.284 0.504 8.356 0.72 ; 
      RECT 8.124 0.504 8.356 0.576 ; 
      RECT 6.86 0.888 7.492 0.96 ; 
      RECT 7.42 0.752 7.492 0.96 ; 
      RECT 7.42 0.752 7.708 0.824 ; 
      RECT 7.636 0.252 7.708 0.824 ; 
      RECT 7.076 0.252 7.708 0.324 ; 
      RECT 5.132 0.892 5.576 0.964 ; 
      RECT 5.504 0.108 5.576 0.964 ; 
      RECT 5.504 0.724 6 0.796 ; 
      RECT 7.42 0.396 7.492 0.588 ; 
      RECT 6.772 0.108 6.844 0.588 ; 
      RECT 6.772 0.396 7.492 0.468 ; 
      RECT 5.348 0.108 6.844 0.18 ; 
      RECT 6.344 0.892 6.544 0.964 ; 
      RECT 6.344 0.308 6.416 0.964 ; 
      RECT 6.344 0.308 6.544 0.38 ; 
      RECT 5.98 0.896 6.196 0.968 ; 
      RECT 6.12 0.292 6.196 0.968 ; 
      RECT 5.676 0.292 6.196 0.364 ; 
      RECT 5.26 0.72 5.404 0.792 ; 
      RECT 5.26 0.288 5.332 0.792 ; 
      RECT 5.136 0.288 5.332 0.36 ; 
      RECT 4.484 0.896 4.9 0.968 ; 
      RECT 4.828 0.108 4.9 0.968 ; 
      RECT 4.464 0.108 4.9 0.18 ; 
      RECT 3.832 0.892 4.032 0.964 ; 
      RECT 3.96 0.308 4.032 0.964 ; 
      RECT 3.832 0.308 4.032 0.38 ; 
      RECT 3.532 0.396 3.604 0.588 ; 
      RECT 2.884 0.396 2.956 0.588 ; 
      RECT 2.884 0.396 3.604 0.468 ; 
      RECT 2.884 0.888 3.516 0.96 ; 
      RECT 2.884 0.752 2.956 0.96 ; 
      RECT 2.668 0.752 2.956 0.824 ; 
      RECT 2.668 0.252 2.74 0.824 ; 
      RECT 2.668 0.252 3.3 0.324 ; 
      RECT 1.676 0.648 2.296 0.72 ; 
      RECT 2.02 0.504 2.092 0.72 ; 
      RECT 2.02 0.504 2.252 0.576 ; 
      RECT 1.652 0.504 1.876 0.576 ; 
      RECT 1.804 0.36 1.876 0.576 ; 
      RECT 1.612 0.36 2.22 0.432 ; 
      RECT 1.372 0.396 1.444 0.588 ; 
      RECT 0.724 0.396 0.796 0.588 ; 
      RECT 0.724 0.396 1.444 0.468 ; 
      RECT 0.724 0.888 1.356 0.96 ; 
      RECT 0.724 0.752 0.796 0.96 ; 
      RECT 0.508 0.752 0.796 0.824 ; 
      RECT 0.508 0.252 0.58 0.824 ; 
      RECT 0.508 0.252 1.14 0.324 ; 
    LAYER M2 ; 
      RECT 1.348 0.432 9.028 0.504 ; 
      RECT 3.932 0.72 6.436 0.792 ; 
    LAYER V1 ; 
      RECT 8.932 0.432 9.004 0.504 ; 
      RECT 6.772 0.432 6.844 0.504 ; 
      RECT 6.344 0.72 6.416 0.792 ; 
      RECT 5.312 0.72 5.384 0.792 ; 
      RECT 3.96 0.72 4.032 0.792 ; 
      RECT 3.532 0.432 3.604 0.504 ; 
      RECT 1.372 0.432 1.444 0.504 ; 
  END 
END ICGx5p33DC_ASAP7_75t_R 


MACRO ICGx6p67DC_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx6p67DC_ASAP7_75t_R 0 0 ; 
  SIZE 10.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 9.864 0.9 10.084 0.972 ; 
        RECT 10.012 0.108 10.084 0.972 ; 
        RECT 9.784 0.108 10.084 0.18 ; 
        RECT 7.704 0.9 7.924 0.972 ; 
        RECT 7.852 0.108 7.924 0.972 ; 
        RECT 7.624 0.108 7.924 0.18 ; 
        RECT 2.452 0.108 2.752 0.18 ; 
        RECT 2.452 0.9 2.672 0.972 ; 
        RECT 2.452 0.108 2.524 0.972 ; 
        RECT 0.292 0.108 0.592 0.18 ; 
        RECT 0.292 0.9 0.512 0.972 ; 
        RECT 0.292 0.108 0.364 0.972 ; 
      LAYER M2 ; 
        RECT 0.248 0.144 10.128 0.216 ; 
      LAYER V1 ; 
        RECT 0.292 0.144 0.364 0.216 ; 
        RECT 2.452 0.144 2.524 0.216 ; 
        RECT 7.852 0.144 7.924 0.216 ; 
        RECT 10.012 0.144 10.084 0.216 ; 
    END 
  END GCLK 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 10.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 10.376 0.036 ; 
    END 
  END VSS 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 9.128 0.684 9.404 0.756 ; 
        RECT 9.332 0.54 9.404 0.756 ; 
        RECT 9.172 0.54 9.404 0.612 ; 
        RECT 6.556 0.712 7.168 0.784 ; 
        RECT 7.096 0.568 7.168 0.784 ; 
        RECT 6.556 0.464 6.628 0.784 ; 
        RECT 5.692 0.576 5.896 0.648 ; 
        RECT 5.692 0.48 5.764 0.648 ; 
        RECT 5.044 0.476 5.116 0.736 ; 
        RECT 3.208 0.712 3.82 0.784 ; 
        RECT 3.748 0.464 3.82 0.784 ; 
        RECT 3.208 0.568 3.28 0.784 ; 
        RECT 0.996 0.684 1.272 0.756 ; 
        RECT 0.996 0.54 1.228 0.612 ; 
        RECT 0.996 0.54 1.068 0.756 ; 
      LAYER M2 ; 
        RECT 0.944 0.576 9.436 0.648 ; 
      LAYER V1 ; 
        RECT 0.996 0.576 1.068 0.648 ; 
        RECT 3.748 0.576 3.82 0.648 ; 
        RECT 5.044 0.576 5.116 0.648 ; 
        RECT 5.764 0.576 5.836 0.648 ; 
        RECT 6.556 0.576 6.628 0.648 ; 
        RECT 9.332 0.576 9.404 0.648 ; 
    END 
  END CLK 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.308 0.688 4.468 0.796 ; 
        RECT 4.396 0.28 4.468 0.796 ; 
        RECT 4.132 0.888 4.384 0.964 ; 
        RECT 4.308 0.688 4.384 0.964 ; 
      LAYER M2 ; 
        RECT 3.932 0.864 4.952 0.936 ; 
      LAYER V1 ; 
        RECT 4.308 0.864 4.384 0.936 ; 
    END 
  END ENA 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.612 0.28 4.684 0.796 ; 
      LAYER M2 ; 
        RECT 3.932 0.288 4.952 0.36 ; 
      LAYER V1 ; 
        RECT 4.612 0.288 4.684 0.36 ; 
    END 
  END SE 
  OBS 
    LAYER M1 ; 
      RECT 9.02 0.888 9.652 0.96 ; 
      RECT 9.58 0.752 9.652 0.96 ; 
      RECT 9.58 0.752 9.868 0.824 ; 
      RECT 9.796 0.252 9.868 0.824 ; 
      RECT 9.236 0.252 9.868 0.324 ; 
      RECT 9.58 0.396 9.652 0.588 ; 
      RECT 8.932 0.396 9.004 0.588 ; 
      RECT 8.932 0.396 9.652 0.468 ; 
      RECT 8.5 0.504 8.724 0.576 ; 
      RECT 8.5 0.36 8.572 0.576 ; 
      RECT 8.156 0.36 8.764 0.432 ; 
      RECT 8.08 0.648 8.7 0.72 ; 
      RECT 8.284 0.504 8.356 0.72 ; 
      RECT 8.124 0.504 8.356 0.576 ; 
      RECT 6.86 0.888 7.492 0.96 ; 
      RECT 7.42 0.752 7.492 0.96 ; 
      RECT 7.42 0.752 7.708 0.824 ; 
      RECT 7.636 0.252 7.708 0.824 ; 
      RECT 7.076 0.252 7.708 0.324 ; 
      RECT 5.132 0.892 5.576 0.964 ; 
      RECT 5.504 0.108 5.576 0.964 ; 
      RECT 5.504 0.724 6 0.796 ; 
      RECT 7.42 0.396 7.492 0.588 ; 
      RECT 6.772 0.108 6.844 0.588 ; 
      RECT 6.772 0.396 7.492 0.468 ; 
      RECT 5.348 0.108 6.844 0.18 ; 
      RECT 6.344 0.892 6.544 0.964 ; 
      RECT 6.344 0.308 6.416 0.964 ; 
      RECT 6.344 0.308 6.544 0.38 ; 
      RECT 5.98 0.896 6.196 0.968 ; 
      RECT 6.12 0.292 6.196 0.968 ; 
      RECT 5.676 0.292 6.196 0.364 ; 
      RECT 5.26 0.72 5.404 0.792 ; 
      RECT 5.26 0.288 5.332 0.792 ; 
      RECT 5.136 0.288 5.332 0.36 ; 
      RECT 4.484 0.896 4.9 0.968 ; 
      RECT 4.828 0.108 4.9 0.968 ; 
      RECT 4.464 0.108 4.9 0.18 ; 
      RECT 3.832 0.892 4.032 0.964 ; 
      RECT 3.96 0.308 4.032 0.964 ; 
      RECT 3.832 0.308 4.032 0.38 ; 
      RECT 3.532 0.396 3.604 0.588 ; 
      RECT 2.884 0.396 2.956 0.588 ; 
      RECT 2.884 0.396 3.604 0.468 ; 
      RECT 2.884 0.888 3.516 0.96 ; 
      RECT 2.884 0.752 2.956 0.96 ; 
      RECT 2.668 0.752 2.956 0.824 ; 
      RECT 2.668 0.252 2.74 0.824 ; 
      RECT 2.668 0.252 3.3 0.324 ; 
      RECT 1.676 0.648 2.296 0.72 ; 
      RECT 2.02 0.504 2.092 0.72 ; 
      RECT 2.02 0.504 2.252 0.576 ; 
      RECT 1.652 0.504 1.876 0.576 ; 
      RECT 1.804 0.36 1.876 0.576 ; 
      RECT 1.612 0.36 2.22 0.432 ; 
      RECT 1.372 0.396 1.444 0.588 ; 
      RECT 0.724 0.396 0.796 0.588 ; 
      RECT 0.724 0.396 1.444 0.468 ; 
      RECT 0.724 0.888 1.356 0.96 ; 
      RECT 0.724 0.752 0.796 0.96 ; 
      RECT 0.508 0.752 0.796 0.824 ; 
      RECT 0.508 0.252 0.58 0.824 ; 
      RECT 0.508 0.252 1.14 0.324 ; 
    LAYER M2 ; 
      RECT 1.348 0.432 9.028 0.504 ; 
      RECT 3.932 0.72 6.436 0.792 ; 
    LAYER V1 ; 
      RECT 8.932 0.432 9.004 0.504 ; 
      RECT 6.772 0.432 6.844 0.504 ; 
      RECT 6.344 0.72 6.416 0.792 ; 
      RECT 5.312 0.72 5.384 0.792 ; 
      RECT 3.96 0.72 4.032 0.792 ; 
      RECT 3.532 0.432 3.604 0.504 ; 
      RECT 1.372 0.432 1.444 0.504 ; 
  END 
END ICGx6p67DC_ASAP7_75t_R 


MACRO ICGx8DC_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN ICGx8DC_ASAP7_75t_R 0 0 ; 
  SIZE 10.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN GCLK 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 9.864 0.9 10.084 0.972 ; 
        RECT 10.012 0.108 10.084 0.972 ; 
        RECT 9.784 0.108 10.084 0.18 ; 
        RECT 7.704 0.9 7.924 0.972 ; 
        RECT 7.852 0.108 7.924 0.972 ; 
        RECT 7.624 0.108 7.924 0.18 ; 
        RECT 2.452 0.108 2.752 0.18 ; 
        RECT 2.452 0.9 2.672 0.972 ; 
        RECT 2.452 0.108 2.524 0.972 ; 
        RECT 0.292 0.108 0.592 0.18 ; 
        RECT 0.292 0.9 0.512 0.972 ; 
        RECT 0.292 0.108 0.364 0.972 ; 
      LAYER M2 ; 
        RECT 0.248 0.144 10.128 0.216 ; 
      LAYER V1 ; 
        RECT 0.292 0.144 0.364 0.216 ; 
        RECT 2.452 0.144 2.524 0.216 ; 
        RECT 7.852 0.144 7.924 0.216 ; 
        RECT 10.012 0.144 10.084 0.216 ; 
    END 
  END GCLK 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 10.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 10.376 0.036 ; 
    END 
  END VSS 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 9.128 0.684 9.404 0.756 ; 
        RECT 9.332 0.54 9.404 0.756 ; 
        RECT 9.172 0.54 9.404 0.612 ; 
        RECT 6.556 0.712 7.168 0.784 ; 
        RECT 7.096 0.568 7.168 0.784 ; 
        RECT 6.556 0.464 6.628 0.784 ; 
        RECT 5.692 0.576 5.896 0.648 ; 
        RECT 5.692 0.48 5.764 0.648 ; 
        RECT 5.044 0.476 5.116 0.736 ; 
        RECT 3.208 0.712 3.82 0.784 ; 
        RECT 3.748 0.464 3.82 0.784 ; 
        RECT 3.208 0.568 3.28 0.784 ; 
        RECT 0.996 0.684 1.272 0.756 ; 
        RECT 0.996 0.54 1.228 0.612 ; 
        RECT 0.996 0.54 1.068 0.756 ; 
      LAYER M2 ; 
        RECT 0.944 0.576 9.436 0.648 ; 
      LAYER V1 ; 
        RECT 0.996 0.576 1.068 0.648 ; 
        RECT 3.748 0.576 3.82 0.648 ; 
        RECT 5.044 0.576 5.116 0.648 ; 
        RECT 5.764 0.576 5.836 0.648 ; 
        RECT 6.556 0.576 6.628 0.648 ; 
        RECT 9.332 0.576 9.404 0.648 ; 
    END 
  END CLK 
  PIN ENA 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.308 0.688 4.468 0.796 ; 
        RECT 4.396 0.28 4.468 0.796 ; 
        RECT 4.132 0.888 4.384 0.964 ; 
        RECT 4.308 0.688 4.384 0.964 ; 
      LAYER M2 ; 
        RECT 3.932 0.864 4.952 0.936 ; 
      LAYER V1 ; 
        RECT 4.308 0.864 4.384 0.936 ; 
    END 
  END ENA 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 4.612 0.28 4.684 0.796 ; 
      LAYER M2 ; 
        RECT 3.932 0.288 4.952 0.36 ; 
      LAYER V1 ; 
        RECT 4.612 0.288 4.684 0.36 ; 
    END 
  END SE 
  OBS 
    LAYER M1 ; 
      RECT 9.02 0.888 9.652 0.96 ; 
      RECT 9.58 0.752 9.652 0.96 ; 
      RECT 9.58 0.752 9.868 0.824 ; 
      RECT 9.796 0.252 9.868 0.824 ; 
      RECT 9.236 0.252 9.868 0.324 ; 
      RECT 9.58 0.396 9.652 0.588 ; 
      RECT 8.932 0.396 9.004 0.588 ; 
      RECT 8.932 0.396 9.652 0.468 ; 
      RECT 8.5 0.504 8.724 0.576 ; 
      RECT 8.5 0.36 8.572 0.576 ; 
      RECT 8.156 0.36 8.764 0.432 ; 
      RECT 8.08 0.648 8.7 0.72 ; 
      RECT 8.284 0.504 8.356 0.72 ; 
      RECT 8.124 0.504 8.356 0.576 ; 
      RECT 6.86 0.888 7.492 0.96 ; 
      RECT 7.42 0.752 7.492 0.96 ; 
      RECT 7.42 0.752 7.708 0.824 ; 
      RECT 7.636 0.252 7.708 0.824 ; 
      RECT 7.076 0.252 7.708 0.324 ; 
      RECT 5.132 0.892 5.576 0.964 ; 
      RECT 5.504 0.108 5.576 0.964 ; 
      RECT 5.504 0.724 6 0.796 ; 
      RECT 7.42 0.396 7.492 0.588 ; 
      RECT 6.772 0.108 6.844 0.588 ; 
      RECT 6.772 0.396 7.492 0.468 ; 
      RECT 5.348 0.108 6.844 0.18 ; 
      RECT 6.344 0.892 6.544 0.964 ; 
      RECT 6.344 0.308 6.416 0.964 ; 
      RECT 6.344 0.308 6.544 0.38 ; 
      RECT 5.98 0.896 6.196 0.968 ; 
      RECT 6.12 0.292 6.196 0.968 ; 
      RECT 5.676 0.292 6.196 0.364 ; 
      RECT 5.26 0.72 5.404 0.792 ; 
      RECT 5.26 0.288 5.332 0.792 ; 
      RECT 5.136 0.288 5.332 0.36 ; 
      RECT 4.484 0.896 4.9 0.968 ; 
      RECT 4.828 0.108 4.9 0.968 ; 
      RECT 4.464 0.108 4.9 0.18 ; 
      RECT 3.832 0.892 4.032 0.964 ; 
      RECT 3.96 0.308 4.032 0.964 ; 
      RECT 3.832 0.308 4.032 0.38 ; 
      RECT 3.532 0.396 3.604 0.588 ; 
      RECT 2.884 0.396 2.956 0.588 ; 
      RECT 2.884 0.396 3.604 0.468 ; 
      RECT 2.884 0.888 3.516 0.96 ; 
      RECT 2.884 0.752 2.956 0.96 ; 
      RECT 2.668 0.752 2.956 0.824 ; 
      RECT 2.668 0.252 2.74 0.824 ; 
      RECT 2.668 0.252 3.3 0.324 ; 
      RECT 1.676 0.648 2.296 0.72 ; 
      RECT 2.02 0.504 2.092 0.72 ; 
      RECT 2.02 0.504 2.252 0.576 ; 
      RECT 1.652 0.504 1.876 0.576 ; 
      RECT 1.804 0.36 1.876 0.576 ; 
      RECT 1.612 0.36 2.22 0.432 ; 
      RECT 1.372 0.396 1.444 0.588 ; 
      RECT 0.724 0.396 0.796 0.588 ; 
      RECT 0.724 0.396 1.444 0.468 ; 
      RECT 0.724 0.888 1.356 0.96 ; 
      RECT 0.724 0.752 0.796 0.96 ; 
      RECT 0.508 0.752 0.796 0.824 ; 
      RECT 0.508 0.252 0.58 0.824 ; 
      RECT 0.508 0.252 1.14 0.324 ; 
    LAYER M2 ; 
      RECT 1.348 0.432 9.028 0.504 ; 
      RECT 3.932 0.72 6.436 0.792 ; 
    LAYER V1 ; 
      RECT 8.932 0.432 9.004 0.504 ; 
      RECT 6.772 0.432 6.844 0.504 ; 
      RECT 6.344 0.72 6.416 0.792 ; 
      RECT 5.312 0.72 5.384 0.792 ; 
      RECT 3.96 0.72 4.032 0.792 ; 
      RECT 3.532 0.432 3.604 0.504 ; 
      RECT 1.372 0.432 1.444 0.504 ; 
  END 
END ICGx8DC_ASAP7_75t_R 


MACRO INVx11_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx11_ASAP7_75t_R 0 0 ; 
  SIZE 2.808 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.808 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.808 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 2.736 0.972 ; 
        RECT 2.664 0.108 2.736 0.972 ; 
        RECT 0.376 0.108 2.736 0.18 ; 
    END 
  END Y 
END INVx11_ASAP7_75t_R 


MACRO INVx13_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx13_ASAP7_75t_R 0 0 ; 
  SIZE 3.24 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.24 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.24 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 3.168 0.972 ; 
        RECT 3.096 0.108 3.168 0.972 ; 
        RECT 0.376 0.108 3.168 0.18 ; 
    END 
  END Y 
END INVx13_ASAP7_75t_R 


MACRO INVx1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx1_ASAP7_75t_R 0 0 ; 
  SIZE 0.648 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.648 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.648 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 0.576 0.972 ; 
        RECT 0.504 0.108 0.576 0.972 ; 
        RECT 0.376 0.108 0.576 0.18 ; 
    END 
  END Y 
END INVx1_ASAP7_75t_R 


MACRO INVx2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx2_ASAP7_75t_R 0 0 ; 
  SIZE 0.864 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.864 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.864 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 0.576 0.972 ; 
        RECT 0.504 0.108 0.576 0.972 ; 
        RECT 0.376 0.108 0.576 0.18 ; 
    END 
  END Y 
END INVx2_ASAP7_75t_R 


MACRO INVx3_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx3_ASAP7_75t_R 0 0 ; 
  SIZE 1.08 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.08 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 1.008 0.972 ; 
        RECT 0.936 0.108 1.008 0.972 ; 
        RECT 0.376 0.108 1.008 0.18 ; 
    END 
  END Y 
END INVx3_ASAP7_75t_R 


MACRO INVx4_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx4_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 1.224 0.972 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
        RECT 0.376 0.108 1.224 0.18 ; 
    END 
  END Y 
END INVx4_ASAP7_75t_R 


MACRO INVx5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx5_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 1.44 0.972 ; 
        RECT 1.368 0.108 1.44 0.972 ; 
        RECT 0.376 0.108 1.44 0.18 ; 
    END 
  END Y 
END INVx5_ASAP7_75t_R 


MACRO INVx6_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx6_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 1.656 0.972 ; 
        RECT 1.584 0.108 1.656 0.972 ; 
        RECT 0.376 0.108 1.656 0.18 ; 
    END 
  END Y 
END INVx6_ASAP7_75t_R 


MACRO INVx8_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVx8_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 2.088 0.972 ; 
        RECT 2.016 0.108 2.088 0.972 ; 
        RECT 0.376 0.108 2.088 0.18 ; 
    END 
  END Y 
END INVx8_ASAP7_75t_R 


MACRO INVxp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVxp33_ASAP7_75t_R 0 0 ; 
  SIZE 0.648 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.136 0.144 0.944 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.648 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.648 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 0.576 0.972 ; 
        RECT 0.504 0.108 0.576 0.972 ; 
        RECT 0.376 0.108 0.576 0.18 ; 
    END 
  END Y 
END INVxp33_ASAP7_75t_R 


MACRO INVxp67_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN INVxp67_ASAP7_75t_R 0 0 ; 
  SIZE 0.648 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.136 0.144 0.944 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.648 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.648 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 0.576 0.972 ; 
        RECT 0.504 0.108 0.576 0.972 ; 
        RECT 0.376 0.108 0.576 0.18 ; 
    END 
  END Y 
END INVxp67_ASAP7_75t_R 


MACRO MAJIxp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MAJIxp5_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.656 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.504 1.028 0.576 ; 
        RECT 0.072 0.756 0.792 0.828 ; 
        RECT 0.72 0.504 0.792 0.828 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.136 0.144 0.828 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.02 0.756 1.444 0.828 ; 
        RECT 1.372 0.252 1.444 0.828 ; 
        RECT 1.02 0.252 1.444 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.108 1.352 0.18 ; 
      RECT 0.376 0.9 1.352 0.972 ; 
  END 
END MAJIxp5_ASAP7_75t_R 


MACRO MAJx2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MAJx2_ASAP7_75t_R 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.424 0.36 0.656 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.756 1.332 0.828 ; 
        RECT 1.26 0.424 1.332 0.828 ; 
        RECT 1.132 0.504 1.332 0.576 ; 
        RECT 0.72 0.504 0.792 0.828 ; 
        RECT 0.484 0.504 0.792 0.576 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.944 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.456 0.9 1.872 0.972 ; 
        RECT 1.8 0.108 1.872 0.972 ; 
        RECT 1.456 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.072 0.756 0.492 0.828 ; 
      RECT 0.072 0.252 0.144 0.828 ; 
      RECT 1.472 0.252 1.544 0.596 ; 
      RECT 0.072 0.252 1.544 0.324 ; 
      RECT 0.16 0.108 1.136 0.18 ; 
      RECT 0.16 0.9 1.136 0.972 ; 
  END 
END MAJx2_ASAP7_75t_R 


MACRO MAJx3_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN MAJx3_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.424 0.36 0.656 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.756 1.332 0.828 ; 
        RECT 1.26 0.424 1.332 0.828 ; 
        RECT 1.132 0.504 1.332 0.576 ; 
        RECT 0.72 0.504 0.792 0.828 ; 
        RECT 0.484 0.504 0.792 0.576 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.456 0.9 2.016 0.972 ; 
        RECT 1.456 0.108 2.016 0.18 ; 
        RECT 1.8 0.108 1.872 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.072 0.756 0.492 0.828 ; 
      RECT 0.072 0.252 0.144 0.828 ; 
      RECT 1.472 0.252 1.544 0.596 ; 
      RECT 0.072 0.252 1.544 0.324 ; 
      RECT 0.16 0.108 1.136 0.18 ; 
      RECT 0.16 0.9 1.136 0.972 ; 
  END 
END MAJx3_ASAP7_75t_R 


MACRO NAND2x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND2x1_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.336 0.576 ; 
        RECT 0.072 0.26 0.144 0.944 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 1.224 0.972 ; 
        RECT 1.152 0.252 1.224 0.972 ; 
        RECT 0.808 0.252 1.224 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 1.136 0.18 ; 
  END 
END NAND2x1_ASAP7_75t_R 


MACRO NAND2x1p5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND2x1p5_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.336 0.576 ; 
        RECT 0.072 0.136 0.144 0.944 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.504 1.028 0.576 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 1.656 0.972 ; 
        RECT 1.584 0.108 1.656 0.972 ; 
        RECT 1.044 0.108 1.656 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.808 0.252 1.352 0.324 ; 
      RECT 0.376 0.108 0.9 0.18 ; 
  END 
END NAND2x1p5_ASAP7_75t_R 


MACRO NAND2x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND2x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.968 0.756 1.116 0.828 ; 
        RECT 1.044 0.424 1.116 0.828 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.396 1.872 0.708 ; 
        RECT 1.288 0.396 1.872 0.468 ; 
        RECT 1.288 0.252 1.36 0.468 ; 
        RECT 0.8 0.252 1.36 0.324 ; 
        RECT 0.288 0.396 0.872 0.468 ; 
        RECT 0.8 0.252 0.872 0.468 ; 
        RECT 0.288 0.756 0.436 0.828 ; 
        RECT 0.288 0.396 0.36 0.828 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 2.088 0.972 ; 
        RECT 2.016 0.252 2.088 0.972 ; 
        RECT 1.672 0.252 2.088 0.324 ; 
        RECT 0.072 0.252 0.488 0.324 ; 
        RECT 0.072 0.252 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 2 0.18 ; 
  END 
END NAND2x2_ASAP7_75t_R 


MACRO NAND2xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND2xp33_ASAP7_75t_R 0 0 ; 
  SIZE 0.864 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.864 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.864 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 0.792 0.972 ; 
        RECT 0.72 0.108 0.792 0.972 ; 
        RECT 0.572 0.108 0.792 0.18 ; 
    END 
  END Y 
END NAND2xp33_ASAP7_75t_R 


MACRO NAND2xp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND2xp5_ASAP7_75t_R 0 0 ; 
  SIZE 0.864 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.424 0.252 0.576 0.324 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.864 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.864 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 0.792 0.972 ; 
        RECT 0.72 0.108 0.792 0.972 ; 
        RECT 0.572 0.108 0.792 0.18 ; 
    END 
  END Y 
END NAND2xp5_ASAP7_75t_R 


MACRO NAND2xp67_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND2xp67_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.5 0.38 0.572 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.252 0.22 0.324 ; 
        RECT 0.072 0.252 0.144 0.972 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.86 0.756 1.008 0.828 ; 
        RECT 0.936 0.424 1.008 0.828 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.9 1.224 0.972 ; 
        RECT 1.152 0.252 1.224 0.972 ; 
        RECT 0.808 0.252 1.224 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 1.136 0.18 ; 
  END 
END NAND2xp67_ASAP7_75t_R 


MACRO NAND3x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND3x1_ASAP7_75t_R 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.608 0.72 1.872 0.792 ; 
        RECT 1.8 0.432 1.872 0.792 ; 
        RECT 1.6 0.432 1.872 0.504 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.972 0.72 1.224 0.792 ; 
        RECT 1.152 0.432 1.224 0.792 ; 
        RECT 0.984 0.432 1.224 0.504 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.244 0.412 0.316 0.812 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.9 2.304 0.972 ; 
        RECT 2.232 0.252 2.304 0.972 ; 
        RECT 1.672 0.252 2.304 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.024 0.108 2 0.18 ; 
      RECT 0.376 0.252 1.352 0.324 ; 
      RECT 0.16 0.108 0.704 0.18 ; 
  END 
END NAND3x1_ASAP7_75t_R 


MACRO NAND3x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND3x2_ASAP7_75t_R 0 0 ; 
  SIZE 4.32 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.352 0.756 2.972 0.828 ; 
        RECT 2.9 0.424 2.972 0.828 ; 
        RECT 1.352 0.424 1.424 0.828 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.188 0.424 2.26 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.32 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.32 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 4.248 0.972 ; 
        RECT 4.176 0.252 4.248 0.972 ; 
        RECT 3.616 0.252 4.248 0.324 ; 
        RECT 0.072 0.252 0.704 0.324 ; 
        RECT 0.072 0.252 0.144 0.972 ; 
    END 
  END Y 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.676 0.72 3.632 0.792 ; 
      LAYER M1 ; 
        RECT 3.464 0.756 3.612 0.828 ; 
        RECT 3.54 0.432 3.612 0.828 ; 
        RECT 0.696 0.756 0.844 0.828 ; 
        RECT 0.696 0.424 0.768 0.828 ; 
      LAYER V1 ; 
        RECT 0.696 0.72 0.768 0.792 ; 
        RECT 3.54 0.72 3.612 0.792 ; 
    END 
  END A 
  OBS 
    LAYER M1 ; 
      RECT 2.968 0.108 3.944 0.18 ; 
      RECT 1.024 0.252 3.296 0.324 ; 
      RECT 1.672 0.108 2.648 0.18 ; 
      RECT 0.376 0.108 1.352 0.18 ; 
  END 
END NAND3x2_ASAP7_75t_R 


MACRO NAND3xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND3xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.08 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.136 0.576 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.136 0.792 0.8 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.08 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.704 0.972 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
END NAND3xp33_ASAP7_75t_R 


MACRO NAND4xp25_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND4xp25_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.136 0.792 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.136 0.576 0.8 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.136 0.36 0.8 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.16 0.9 1.224 0.972 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
        RECT 1.024 0.108 1.224 0.18 ; 
    END 
  END Y 
END NAND4xp25_ASAP7_75t_R 


MACRO NAND4xp75_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND4xp75_ASAP7_75t_R 0 0 ; 
  SIZE 3.024 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.448 0.424 2.52 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.404 2.196 0.476 ; 
        RECT 2.124 0.28 2.196 0.476 ; 
        RECT 2.016 0.404 2.088 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.404 1.224 0.8 ; 
        RECT 0.828 0.404 1.224 0.476 ; 
        RECT 0.828 0.28 0.9 0.476 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.9 0.228 0.972 ; 
        RECT 0.072 0.108 0.228 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.024 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 2.952 0.972 ; 
        RECT 2.88 0.252 2.952 0.972 ; 
        RECT 2.32 0.252 2.952 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.648 0.108 2.664 0.18 ; 
      RECT 1.024 0.252 1.996 0.324 ; 
      RECT 0.368 0.108 1.36 0.18 ; 
  END 
END NAND4xp75_ASAP7_75t_R 


MACRO NAND5xp2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NAND5xp2_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.136 0.576 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.136 0.792 0.8 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.136 1.008 0.8 ; 
    END 
  END D 
  PIN E 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.136 1.224 0.8 ; 
    END 
  END E 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.036 0.9 1.268 0.972 ; 
        RECT 0.036 0.108 0.28 0.18 ; 
        RECT 0.036 0.108 0.108 0.972 ; 
    END 
  END Y 
END NAND5xp2_ASAP7_75t_R 


MACRO NOR2x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR2x1_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.336 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.828 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.504 0.92 0.576 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.756 1.224 0.828 ; 
        RECT 1.152 0.108 1.224 0.828 ; 
        RECT 0.376 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 1.136 0.972 ; 
  END 
END NOR2x1_ASAP7_75t_R 


MACRO NOR2x1p5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR2x1p5_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.336 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.504 1.028 0.576 ; 
        RECT 0.504 0.252 0.652 0.324 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.9 1.656 0.972 ; 
        RECT 1.584 0.108 1.656 0.972 ; 
        RECT 0.376 0.108 1.656 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.808 0.756 1.352 0.828 ; 
      RECT 0.376 0.9 0.9 0.972 ; 
  END 
END NOR2x1p5_ASAP7_75t_R 


MACRO NOR2x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR2x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.252 1.116 0.656 ; 
        RECT 0.968 0.252 1.116 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.288 0.612 1.872 0.684 ; 
        RECT 1.8 0.372 1.872 0.684 ; 
        RECT 0.8 0.756 1.36 0.828 ; 
        RECT 1.288 0.612 1.36 0.828 ; 
        RECT 0.8 0.612 0.872 0.828 ; 
        RECT 0.288 0.612 0.872 0.684 ; 
        RECT 0.288 0.252 0.436 0.324 ; 
        RECT 0.288 0.252 0.36 0.684 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.756 2.088 0.828 ; 
        RECT 2.016 0.108 2.088 0.828 ; 
        RECT 0.072 0.108 2.088 0.18 ; 
        RECT 0.072 0.756 0.488 0.828 ; 
        RECT 0.072 0.108 0.144 0.828 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 2 0.972 ; 
  END 
END NOR2x2_ASAP7_75t_R 


MACRO NOR2xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR2xp33_ASAP7_75t_R 0 0 ; 
  SIZE 0.864 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.9 0.22 0.972 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.864 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.864 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.572 0.9 0.792 0.972 ; 
        RECT 0.72 0.108 0.792 0.972 ; 
        RECT 0.376 0.108 0.792 0.18 ; 
    END 
  END Y 
END NOR2xp33_ASAP7_75t_R 


MACRO NOR2xp67_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR2xp67_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.508 0.38 0.58 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.828 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.504 1.028 0.576 ; 
        RECT 0.504 0.252 0.652 0.324 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.756 1.224 0.828 ; 
        RECT 1.152 0.108 1.224 0.828 ; 
        RECT 0.592 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 1.136 0.972 ; 
  END 
END NOR2xp67_ASAP7_75t_R 


MACRO NOR3x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR3x1_ASAP7_75t_R 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.612 1.872 0.684 ; 
        RECT 1.8 0.252 1.872 0.684 ; 
        RECT 1.584 0.252 1.872 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.612 1.224 0.684 ; 
        RECT 1.152 0.252 1.224 0.684 ; 
        RECT 0.936 0.252 1.224 0.324 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.36 0.576 ; 
        RECT 0.072 0.756 0.22 0.828 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.828 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.672 0.756 2.304 0.828 ; 
        RECT 2.232 0.108 2.304 0.828 ; 
        RECT 0.808 0.108 2.304 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.024 0.9 2 0.972 ; 
      RECT 0.376 0.756 1.352 0.828 ; 
      RECT 0.16 0.9 0.704 0.972 ; 
  END 
END NOR3x1_ASAP7_75t_R 


MACRO NOR3x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR3x2_ASAP7_75t_R 0 0 ; 
  SIZE 4.32 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.9 0.252 2.972 0.656 ; 
        RECT 1.352 0.252 2.972 0.324 ; 
        RECT 1.352 0.252 1.424 0.656 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.188 0.424 2.26 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 4.32 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 4.32 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 3.616 0.756 4.248 0.828 ; 
        RECT 4.176 0.108 4.248 0.828 ; 
        RECT 0.072 0.108 4.248 0.18 ; 
        RECT 0.072 0.756 0.704 0.828 ; 
        RECT 0.072 0.108 0.144 0.828 ; 
    END 
  END Y 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.676 0.288 3.632 0.36 ; 
      LAYER M1 ; 
        RECT 3.54 0.252 3.612 0.648 ; 
        RECT 3.464 0.252 3.612 0.324 ; 
        RECT 0.696 0.252 0.844 0.324 ; 
        RECT 0.696 0.252 0.768 0.656 ; 
      LAYER V1 ; 
        RECT 0.696 0.288 0.768 0.36 ; 
        RECT 3.54 0.288 3.612 0.36 ; 
    END 
  END A 
  OBS 
    LAYER M1 ; 
      RECT 2.968 0.9 3.944 0.972 ; 
      RECT 1.024 0.756 3.296 0.828 ; 
      RECT 1.672 0.9 2.648 0.972 ; 
      RECT 0.376 0.9 1.352 0.972 ; 
  END 
END NOR3x2_ASAP7_75t_R 


MACRO NOR3xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR3xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.08 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.944 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.944 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.08 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.704 0.18 ; 
        RECT 0.072 0.9 0.272 0.972 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
END NOR3xp33_ASAP7_75t_R 


MACRO NOR4xp25_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR4xp25_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.944 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.944 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.944 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.9 1.224 0.972 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
        RECT 0.16 0.108 1.224 0.18 ; 
    END 
  END Y 
END NOR4xp25_ASAP7_75t_R 


MACRO NOR4xp75_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR4xp75_ASAP7_75t_R 0 0 ; 
  SIZE 3.024 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.448 0.28 2.52 0.656 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.124 0.604 2.196 0.8 ; 
        RECT 2.016 0.604 2.196 0.676 ; 
        RECT 2.016 0.28 2.088 0.676 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.604 1.224 0.676 ; 
        RECT 1.152 0.28 1.224 0.676 ; 
        RECT 0.828 0.604 0.9 0.8 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.9 0.228 0.972 ; 
        RECT 0.072 0.108 0.228 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.024 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.024 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.32 0.756 2.952 0.828 ; 
        RECT 2.88 0.108 2.952 0.828 ; 
        RECT 0.376 0.108 2.952 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.648 0.9 2.664 0.972 ; 
      RECT 1.024 0.756 1.996 0.828 ; 
      RECT 0.368 0.9 1.36 0.972 ; 
  END 
END NOR4xp75_ASAP7_75t_R 


MACRO NOR5xp2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN NOR5xp2_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.792 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.944 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.944 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.944 ; 
    END 
  END D 
  PIN E 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.944 ; 
    END 
  END E 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.068 0.108 1.352 0.18 ; 
        RECT 0.068 0.9 0.28 0.972 ; 
        RECT 0.068 0.108 0.148 0.972 ; 
    END 
  END Y 
END NOR5xp2_ASAP7_75t_R 


MACRO O2A1O1Ixp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN O2A1O1Ixp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.424 0.36 0.8 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.824 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.9 1.224 0.972 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
        RECT 0.376 0.108 1.224 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.9 0.972 ; 
      RECT 0.16 0.252 0.704 0.324 ; 
  END 
END O2A1O1Ixp33_ASAP7_75t_R 


MACRO O2A1O1Ixp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN O2A1O1Ixp5_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.252 1.008 0.656 ; 
        RECT 0.288 0.252 1.008 0.324 ; 
        RECT 0.288 0.252 0.36 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.656 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.656 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.456 0.9 1.656 0.972 ; 
        RECT 1.584 0.108 1.656 0.972 ; 
        RECT 1.26 0.108 1.656 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.504 0.756 1.352 0.828 ; 
      RECT 0.592 0.108 1.116 0.18 ; 
      RECT 0.376 0.9 0.92 0.972 ; 
  END 
END O2A1O1Ixp5_ASAP7_75t_R 


MACRO OA211x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA211x2_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.36 0.576 ; 
        RECT 0.072 0.28 0.144 0.8 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.656 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.184 0.9 1.656 0.972 ; 
        RECT 1.584 0.108 1.656 0.972 ; 
        RECT 1.144 0.108 1.656 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 1.008 0.972 ; 
      RECT 0.936 0.756 1.008 0.972 ; 
      RECT 0.936 0.756 1.224 0.828 ; 
      RECT 1.152 0.252 1.224 0.828 ; 
      RECT 0.396 0.252 1.224 0.324 ; 
      RECT 0.16 0.108 0.704 0.18 ; 
  END 
END OA211x2_ASAP7_75t_R 


MACRO OA21x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA21x2_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.28 0.144 0.944 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.8 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.612 0.956 0.684 ; 
        RECT 0.72 0.424 0.792 0.684 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.9 1.44 0.972 ; 
        RECT 1.368 0.108 1.44 0.972 ; 
        RECT 1.024 0.108 1.44 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.592 0.9 0.896 0.972 ; 
      RECT 0.824 0.756 0.896 0.972 ; 
      RECT 0.824 0.756 1.224 0.828 ; 
      RECT 1.152 0.252 1.224 0.828 ; 
      RECT 0.396 0.252 1.224 0.324 ; 
      RECT 0.16 0.108 0.704 0.18 ; 
  END 
END OA21x2_ASAP7_75t_R 


MACRO OA221x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA221x2_ASAP7_75t_R 0 0 ; 
  SIZE 3.456 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.86 0.756 1.008 0.828 ; 
        RECT 0.936 0.396 1.008 0.828 ; 
        RECT 0.86 0.396 1.008 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.756 1.516 0.828 ; 
        RECT 1.368 0.396 1.516 0.468 ; 
        RECT 1.368 0.396 1.44 0.828 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.372 0.756 2.52 0.828 ; 
        RECT 2.448 0.396 2.52 0.828 ; 
        RECT 2.372 0.396 2.52 0.468 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.94 0.756 2.088 0.828 ; 
        RECT 2.016 0.396 2.088 0.828 ; 
        RECT 1.94 0.396 2.088 0.468 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.88 0.756 3.028 0.828 ; 
        RECT 2.88 0.396 3.028 0.468 ; 
        RECT 2.88 0.396 2.952 0.828 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.456 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.456 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.488 0.18 ; 
        RECT 0.072 0.9 0.468 0.972 ; 
        RECT 0.396 0.756 0.468 0.972 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.576 0.9 3.384 0.972 ; 
      RECT 3.312 0.252 3.384 0.972 ; 
      RECT 0.576 0.504 0.648 0.972 ; 
      RECT 0.484 0.504 0.648 0.576 ; 
      RECT 2.964 0.252 3.384 0.324 ; 
      RECT 1.888 0.108 3.296 0.18 ; 
      RECT 0.808 0.252 2.672 0.324 ; 
  END 
END OA221x2_ASAP7_75t_R 


MACRO OA222x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA222x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.424 0.36 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.8 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.8 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.28 1.872 0.8 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.592 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.124 0.9 2.52 0.972 ; 
        RECT 2.448 0.108 2.52 0.972 ; 
        RECT 2.104 0.108 2.52 0.18 ; 
        RECT 2.124 0.756 2.196 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.036 0.9 2.016 0.972 ; 
      RECT 1.944 0.504 2.016 0.972 ; 
      RECT 0.036 0.252 0.108 0.972 ; 
      RECT 1.944 0.504 2.216 0.576 ; 
      RECT 0.036 0.252 0.488 0.324 ; 
      RECT 0.808 0.252 1.44 0.324 ; 
      RECT 1.368 0.108 1.44 0.324 ; 
      RECT 1.368 0.108 1.872 0.18 ; 
      RECT 0.16 0.108 1.136 0.18 ; 
  END 
END OA222x2_ASAP7_75t_R 


MACRO OA22x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA22x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.424 1.44 0.8 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.28 1.872 0.944 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.252 1.656 0.8 ; 
        RECT 1.468 0.252 1.656 0.324 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.284 0.9 0.488 0.972 ; 
        RECT 0.284 0.108 0.488 0.18 ; 
        RECT 0.284 0.108 0.364 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.72 0.9 1.568 0.972 ; 
      RECT 0.72 0.252 0.792 0.972 ; 
      RECT 0.548 0.504 0.792 0.576 ; 
      RECT 0.72 0.252 1.332 0.324 ; 
      RECT 1.024 0.108 2 0.18 ; 
  END 
END OA22x2_ASAP7_75t_R 


MACRO OA31x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA31x2_ASAP7_75t_R 0 0 ; 
  SIZE 3.24 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.212 0.756 0.36 0.828 ; 
        RECT 0.288 0.396 0.36 0.828 ; 
        RECT 0.212 0.396 0.36 0.468 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.504 0.812 0.576 ; 
        RECT 0.504 0.756 0.652 0.828 ; 
        RECT 0.504 0.424 0.576 0.828 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.504 1.656 0.576 ; 
        RECT 1.368 0.252 1.44 0.656 ; 
        RECT 1.292 0.252 1.44 0.324 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.94 0.612 2.088 0.684 ; 
        RECT 2.016 0.424 2.088 0.684 ; 
    END 
  END B1 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 3.24 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 3.24 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.772 0.9 3.168 0.972 ; 
        RECT 3.096 0.108 3.168 0.972 ; 
        RECT 2.772 0.108 3.168 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.476 0.756 2.304 0.828 ; 
      RECT 2.232 0.252 2.304 0.828 ; 
      RECT 2.232 0.504 2.668 0.576 ; 
      RECT 1.672 0.252 2.304 0.324 ; 
      RECT 1.268 0.9 1.784 0.972 ; 
      RECT 1.268 0.756 1.34 0.972 ; 
      RECT 0.808 0.756 1.34 0.828 ; 
      RECT 0.376 0.108 2 0.18 ; 
      RECT 0.16 0.252 1.136 0.324 ; 
      RECT 0.16 0.9 1.136 0.972 ; 
  END 
END OA31x2_ASAP7_75t_R 


MACRO OA331x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA331x1_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.664 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.424 1.44 0.8 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.424 1.656 0.8 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.424 1.872 0.8 ; 
    END 
  END C1 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.272 0.972 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.9 2.088 0.972 ; 
      RECT 2.016 0.252 2.088 0.972 ; 
      RECT 0.396 0.744 0.468 0.972 ; 
      RECT 0.288 0.744 0.468 0.816 ; 
      RECT 0.288 0.46 0.36 0.816 ; 
      RECT 1.884 0.252 2.088 0.324 ; 
      RECT 0.936 0.252 1.572 0.324 ; 
      RECT 0.936 0.108 1.008 0.324 ; 
      RECT 0.592 0.108 1.008 0.18 ; 
      RECT 1.232 0.108 1.788 0.18 ; 
  END 
END OA331x1_ASAP7_75t_R 


MACRO OA331x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA331x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.664 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.424 1.44 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.424 1.656 0.8 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.424 1.872 0.8 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.424 2.088 0.8 ; 
    END 
  END C1 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.18 0.9 0.488 0.972 ; 
        RECT 0.18 0.108 0.488 0.18 ; 
        RECT 0.18 0.108 0.252 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.612 0.9 2.304 0.972 ; 
      RECT 2.232 0.252 2.304 0.972 ; 
      RECT 0.612 0.744 0.684 0.972 ; 
      RECT 0.504 0.744 0.684 0.816 ; 
      RECT 0.504 0.46 0.576 0.816 ; 
      RECT 2.1 0.252 2.304 0.324 ; 
      RECT 1.152 0.252 1.788 0.324 ; 
      RECT 1.152 0.108 1.224 0.324 ; 
      RECT 0.808 0.108 1.224 0.18 ; 
      RECT 1.448 0.108 2.004 0.18 ; 
  END 
END OA331x2_ASAP7_75t_R 


MACRO OA332x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA332x1_ASAP7_75t_R 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.656 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.424 1.44 0.8 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.424 1.656 0.8 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.424 2.088 0.8 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.424 1.872 0.8 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.376 0.972 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.504 0.9 2.304 0.972 ; 
      RECT 2.232 0.252 2.304 0.972 ; 
      RECT 0.504 0.756 0.576 0.972 ; 
      RECT 0.288 0.756 0.576 0.828 ; 
      RECT 0.288 0.476 0.36 0.828 ; 
      RECT 1.884 0.252 2.304 0.324 ; 
      RECT 0.936 0.252 1.572 0.324 ; 
      RECT 0.936 0.108 1.008 0.324 ; 
      RECT 0.584 0.108 1.008 0.18 ; 
      RECT 1.232 0.108 2.224 0.18 ; 
  END 
END OA332x1_ASAP7_75t_R 


MACRO OA332x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA332x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.424 1.44 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.424 1.656 0.8 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.424 1.872 0.8 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.232 0.424 2.304 0.8 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.424 2.088 0.8 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.592 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.548 0.972 ; 
        RECT 0.072 0.108 0.488 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.72 0.9 2.52 0.972 ; 
      RECT 2.448 0.252 2.52 0.972 ; 
      RECT 0.72 0.756 0.792 0.972 ; 
      RECT 0.504 0.756 0.792 0.828 ; 
      RECT 0.504 0.476 0.576 0.828 ; 
      RECT 2.1 0.252 2.52 0.324 ; 
      RECT 1.152 0.252 1.788 0.324 ; 
      RECT 1.152 0.108 1.224 0.324 ; 
      RECT 0.8 0.108 1.224 0.18 ; 
      RECT 1.448 0.108 2.44 0.18 ; 
  END 
END OA332x2_ASAP7_75t_R 


MACRO OA333x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA333x1_ASAP7_75t_R 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.232 0.424 2.304 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.424 2.088 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.424 1.872 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.424 1.44 0.8 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.424 1.656 0.8 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END C2 
  PIN C3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.656 ; 
    END 
  END C3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.592 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.272 0.972 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.9 2.52 0.972 ; 
      RECT 2.448 0.252 2.52 0.972 ; 
      RECT 0.396 0.744 0.468 0.972 ; 
      RECT 0.288 0.744 0.468 0.816 ; 
      RECT 0.288 0.46 0.36 0.816 ; 
      RECT 1.868 0.252 2.52 0.324 ; 
      RECT 0.928 0.252 1.576 0.324 ; 
      RECT 0.928 0.108 1 0.324 ; 
      RECT 0.588 0.108 1 0.18 ; 
      RECT 1.236 0.108 2.276 0.18 ; 
  END 
END OA333x1_ASAP7_75t_R 


MACRO OA333x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA333x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.808 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.448 0.424 2.52 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.232 0.424 2.304 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.424 2.088 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.424 1.44 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.424 1.656 0.8 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.424 1.872 0.8 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.8 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END C2 
  PIN C3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.656 ; 
    END 
  END C3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.808 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.808 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.9 0.488 0.972 ; 
        RECT 0.288 0.108 0.488 0.18 ; 
        RECT 0.288 0.108 0.36 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.612 0.9 2.736 0.972 ; 
      RECT 2.664 0.252 2.736 0.972 ; 
      RECT 0.612 0.744 0.684 0.972 ; 
      RECT 0.504 0.744 0.684 0.816 ; 
      RECT 0.504 0.46 0.576 0.816 ; 
      RECT 2.084 0.252 2.736 0.324 ; 
      RECT 1.144 0.252 1.792 0.324 ; 
      RECT 1.144 0.108 1.216 0.324 ; 
      RECT 0.804 0.108 1.216 0.18 ; 
      RECT 1.452 0.108 2.492 0.18 ; 
  END 
END OA333x2_ASAP7_75t_R 


MACRO OA33x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OA33x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.424 1.872 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.424 1.656 0.8 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.424 1.44 0.8 ; 
    END 
  END B3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.108 0.488 0.18 ; 
        RECT 0.072 0.9 0.468 0.972 ; 
        RECT 0.396 0.756 0.468 0.972 ; 
        RECT 0.248 0.756 0.468 0.828 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.576 0.9 2.088 0.972 ; 
      RECT 2.016 0.252 2.088 0.972 ; 
      RECT 0.576 0.504 0.648 0.972 ; 
      RECT 0.484 0.504 0.648 0.576 ; 
      RECT 1.456 0.252 2.088 0.324 ; 
      RECT 0.808 0.108 1.784 0.18 ; 
  END 
END OA33x2_ASAP7_75t_R 


MACRO OAI211xp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI211xp5_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.36 0.576 ; 
        RECT 0.072 0.28 0.144 0.8 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.16 0.9 1.224 0.972 ; 
        RECT 1.152 0.252 1.224 0.972 ; 
        RECT 0.396 0.252 1.224 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 0.704 0.18 ; 
  END 
END OAI211xp5_ASAP7_75t_R 


MACRO OAI21x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21x1_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.756 1.224 0.828 ; 
        RECT 1.152 0.424 1.224 0.828 ; 
        RECT 0.504 0.424 0.576 0.828 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.76 0.508 1.024 0.58 ; 
        RECT 0.76 0.396 0.908 0.684 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.252 1.44 0.616 ; 
        RECT 0.288 0.252 1.44 0.324 ; 
        RECT 0.288 0.252 0.36 0.8 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 1.656 0.972 ; 
        RECT 1.584 0.108 1.656 0.972 ; 
        RECT 1.476 0.108 1.656 0.18 ; 
        RECT 0.072 0.108 0.252 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.108 1.332 0.18 ; 
  END 
END OAI21x1_ASAP7_75t_R 


MACRO OAI21xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.08 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.28 0.144 0.944 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.812 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.08 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.9 1.008 0.972 ; 
        RECT 0.936 0.252 1.008 0.972 ; 
        RECT 0.396 0.252 1.008 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 0.704 0.18 ; 
  END 
END OAI21xp33_ASAP7_75t_R 


MACRO OAI21xp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI21xp5_ASAP7_75t_R 0 0 ; 
  SIZE 1.08 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.28 0.144 0.944 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.812 ; 
    END 
  END A2 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.684 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.08 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.08 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.592 0.9 1.008 0.972 ; 
        RECT 0.936 0.252 1.008 0.972 ; 
        RECT 0.396 0.252 1.008 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 0.704 0.18 ; 
  END 
END OAI21xp5_ASAP7_75t_R 


MACRO OAI221xp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI221xp5_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.944 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.424 0.36 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.8 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.92 0.972 ; 
        RECT 0.072 0.252 0.492 0.324 ; 
        RECT 0.072 0.252 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.804 0.252 1.356 0.324 ; 
      RECT 0.16 0.108 0.704 0.18 ; 
  END 
END OAI221xp5_ASAP7_75t_R 


MACRO OAI222xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI222xp33_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.424 0.36 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.8 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.28 1.656 0.8 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.28 1.872 0.8 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 2.088 0.972 ; 
        RECT 2.016 0.22 2.088 0.972 ; 
        RECT 0.072 0.252 0.488 0.324 ; 
        RECT 0.072 0.252 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.808 0.252 1.44 0.324 ; 
      RECT 1.368 0.108 1.44 0.324 ; 
      RECT 1.368 0.108 1.872 0.18 ; 
      RECT 0.16 0.108 1.136 0.18 ; 
  END 
END OAI222xp33_ASAP7_75t_R 


MACRO OAI22x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI22x1_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.612 1.516 0.684 ; 
        RECT 1.368 0.396 1.516 0.468 ; 
        RECT 1.368 0.396 1.44 0.684 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.756 1.872 0.828 ; 
        RECT 1.8 0.396 1.872 0.828 ; 
        RECT 1.724 0.396 1.872 0.468 ; 
        RECT 1.152 0.472 1.224 0.828 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.644 0.612 0.792 0.684 ; 
        RECT 0.72 0.252 0.792 0.684 ; 
        RECT 0.644 0.252 0.792 0.324 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.756 1.008 0.828 ; 
        RECT 0.936 0.464 1.008 0.828 ; 
        RECT 0.288 0.252 0.436 0.324 ; 
        RECT 0.288 0.252 0.36 0.828 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.152 0.9 2.088 0.972 ; 
        RECT 2.016 0.252 2.088 0.972 ; 
        RECT 1.236 0.252 2.088 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 2 0.18 ; 
  END 
END OAI22x1_ASAP7_75t_R 


MACRO OAI22xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI22xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.424 0.36 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.8 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.9 1.1 0.972 ; 
        RECT 0.936 0.28 1.008 0.972 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.704 0.972 ; 
        RECT 0.072 0.252 0.468 0.324 ; 
        RECT 0.072 0.252 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 1.136 0.18 ; 
  END 
END OAI22xp33_ASAP7_75t_R 


MACRO OAI22xp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI22xp5_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.424 0.36 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.8 ; 
    END 
  END A2 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.9 1.1 0.972 ; 
        RECT 0.936 0.28 1.008 0.972 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.252 0.792 0.656 ; 
        RECT 0.604 0.252 0.792 0.324 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.704 0.972 ; 
        RECT 0.072 0.252 0.468 0.324 ; 
        RECT 0.072 0.252 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.108 1.136 0.18 ; 
  END 
END OAI22xp5_ASAP7_75t_R 


MACRO OAI311xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI311xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.944 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.136 0.144 0.944 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.8 ; 
    END 
  END B1 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.8 ; 
    END 
  END C1 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.792 0.9 1.44 0.972 ; 
        RECT 1.368 0.108 1.44 0.972 ; 
        RECT 1.24 0.108 1.44 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.108 0.936 0.18 ; 
  END 
END OAI311xp33_ASAP7_75t_R 


MACRO OAI31xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI31xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.944 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.944 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.804 0.9 1.224 0.972 ; 
        RECT 1.152 0.252 1.224 0.972 ; 
        RECT 1.024 0.252 1.224 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.372 0.108 0.92 0.18 ; 
  END 
END OAI31xp33_ASAP7_75t_R 


MACRO OAI31xp67_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI31xp67_ASAP7_75t_R 0 0 ; 
  SIZE 2.808 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.664 0.504 2.736 0.792 ; 
        RECT 2.212 0.504 2.736 0.576 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.504 1.676 0.576 ; 
        RECT 1.152 0.504 1.224 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.28 0.144 0.944 ; 
    END 
  END A3 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.504 0.812 0.576 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.808 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.808 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.808 0.252 2.652 0.324 ; 
        RECT 0.808 0.756 1.008 0.828 ; 
        RECT 0.936 0.252 1.008 0.828 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 2.104 0.9 2.652 0.972 ; 
      RECT 1.456 0.756 2.432 0.828 ; 
      RECT 0.16 0.108 2.216 0.18 ; 
      RECT 0.376 0.9 1.784 0.972 ; 
  END 
END OAI31xp67_ASAP7_75t_R 


MACRO OAI321xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI321xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.944 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.38 0.576 ; 
        RECT 0.072 0.136 0.144 0.944 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.424 1.44 0.8 ; 
    END 
  END B2 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.792 0.9 1.656 0.972 ; 
        RECT 1.584 0.252 1.656 0.972 ; 
        RECT 1.24 0.252 1.656 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.024 0.108 1.584 0.18 ; 
      RECT 0.376 0.252 0.92 0.324 ; 
  END 
END OAI321xp33_ASAP7_75t_R 


MACRO OAI322xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI322xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.42 1.224 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.424 0.36 0.944 ; 
    END 
  END B2 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.424 1.656 0.8 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.42 1.44 0.8 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.944 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.588 0.9 1.872 0.972 ; 
        RECT 1.8 0.252 1.872 0.972 ; 
        RECT 1.456 0.252 1.872 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.808 0.108 1.8 0.18 ; 
      RECT 0.156 0.252 1.136 0.324 ; 
  END 
END OAI322xp33_ASAP7_75t_R 


MACRO OAI32xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI32xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.252 0.888 0.324 ; 
        RECT 0.72 0.252 0.792 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.8 ; 
    END 
  END B2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.16 0.9 1.44 0.972 ; 
        RECT 1.368 0.252 1.44 0.972 ; 
        RECT 1.024 0.252 1.44 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.396 0.108 1.352 0.18 ; 
  END 
END OAI32xp33_ASAP7_75t_R 


MACRO OAI331xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI331xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.944 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.424 0.36 0.944 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.8 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.424 1.44 0.8 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.424 1.656 0.8 ; 
    END 
  END C1 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.944 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.804 0.9 1.872 0.972 ; 
        RECT 1.8 0.252 1.872 0.972 ; 
        RECT 1.668 0.252 1.872 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.016 0.108 1.572 0.18 ; 
      RECT 0.368 0.252 1.356 0.324 ; 
  END 
END OAI331xp33_ASAP7_75t_R 


MACRO OAI332xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI332xp33_ASAP7_75t_R 0 0 ; 
  SIZE 2.16 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.944 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.424 0.36 0.944 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.8 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.424 1.44 0.8 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.424 1.872 0.8 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.424 1.656 0.8 ; 
    END 
  END C2 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.16 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.16 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.804 0.9 2.088 0.972 ; 
        RECT 2.016 0.252 2.088 0.972 ; 
        RECT 1.668 0.252 2.088 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.016 0.108 2.008 0.18 ; 
      RECT 0.368 0.252 1.356 0.324 ; 
  END 
END OAI332xp33_ASAP7_75t_R 


MACRO OAI333xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI333xp33_ASAP7_75t_R 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.016 0.424 2.088 0.8 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.424 1.872 0.8 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.424 1.656 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.8 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.424 1.44 0.8 ; 
    END 
  END B3 
  PIN C1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.8 ; 
    END 
  END C1 
  PIN C2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.944 ; 
    END 
  END C2 
  PIN C3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.424 0.36 0.944 ; 
    END 
  END C3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.804 0.9 2.304 0.972 ; 
        RECT 2.232 0.252 2.304 0.972 ; 
        RECT 1.652 0.252 2.304 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.016 0.108 2.06 0.18 ; 
      RECT 0.376 0.252 1.36 0.324 ; 
  END 
END OAI333xp33_ASAP7_75t_R 


MACRO OAI33xp33_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OAI33xp33_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.944 ; 
    END 
  END A1 
  PIN A2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.944 ; 
    END 
  END A2 
  PIN A3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END A3 
  PIN B1 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.424 1.008 0.8 ; 
    END 
  END B1 
  PIN B2 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.8 ; 
    END 
  END B2 
  PIN B3 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.424 1.44 0.8 ; 
    END 
  END B3 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.804 0.9 1.656 0.972 ; 
        RECT 1.584 0.252 1.656 0.972 ; 
        RECT 1.024 0.252 1.656 0.324 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.368 0.108 1.352 0.18 ; 
  END 
END OAI33xp33_ASAP7_75t_R 


MACRO OR2x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x2_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.308 0.576 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.8 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.9 1.224 0.972 ; 
        RECT 1.152 0.108 1.224 0.972 ; 
        RECT 0.828 0.108 1.224 0.18 ; 
        RECT 0.828 0.736 0.9 0.972 ; 
        RECT 0.828 0.108 0.9 0.344 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.744 0.972 ; 
      RECT 0.672 0.108 0.744 0.972 ; 
      RECT 0.672 0.504 0.908 0.576 ; 
      RECT 0.376 0.108 0.744 0.18 ; 
  END 
END OR2x2_ASAP7_75t_R 


MACRO OR2x4_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x4_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.504 0.308 0.576 ; 
        RECT 0.072 0.108 0.22 0.18 ; 
        RECT 0.072 0.108 0.144 0.8 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.9 1.656 0.972 ; 
        RECT 1.584 0.108 1.656 0.972 ; 
        RECT 0.828 0.108 1.656 0.18 ; 
        RECT 1.26 0.736 1.332 0.972 ; 
        RECT 1.26 0.108 1.332 0.344 ; 
        RECT 0.828 0.736 0.9 0.972 ; 
        RECT 0.828 0.108 0.9 0.344 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.748 0.972 ; 
      RECT 0.676 0.108 0.748 0.972 ; 
      RECT 0.676 0.504 0.908 0.576 ; 
      RECT 0.376 0.108 0.748 0.18 ; 
  END 
END OR2x4_ASAP7_75t_R 


MACRO OR2x6_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR2x6_ASAP7_75t_R 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.252 0.576 0.488 ; 
        RECT 0.072 0.252 0.576 0.324 ; 
        RECT 0.072 0.252 0.144 0.944 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.612 1.008 0.684 ; 
        RECT 0.936 0.484 1.008 0.684 ; 
        RECT 0.288 0.424 0.36 0.944 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.592 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.9 2.52 0.972 ; 
        RECT 2.448 0.108 2.52 0.972 ; 
        RECT 1.24 0.108 2.52 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.592 0.756 1.224 0.828 ; 
      RECT 1.152 0.28 1.224 0.828 ; 
      RECT 0.936 0.28 1.224 0.352 ; 
      RECT 0.936 0.108 1.008 0.352 ; 
      RECT 0.376 0.108 1.008 0.18 ; 
  END 
END OR2x6_ASAP7_75t_R 


MACRO OR3x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR3x1_ASAP7_75t_R 0 0 ; 
  SIZE 1.296 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.296 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.296 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.732 1.224 0.804 ; 
        RECT 1.152 0.304 1.224 0.804 ; 
        RECT 1.044 0.304 1.224 0.376 ; 
        RECT 1.044 0.732 1.116 0.94 ; 
        RECT 1.044 0.136 1.116 0.376 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.936 0.972 ; 
      RECT 0.864 0.108 0.936 0.972 ; 
      RECT 0.864 0.504 1.048 0.576 ; 
      RECT 0.16 0.108 0.936 0.18 ; 
  END 
END OR3x1_ASAP7_75t_R 


MACRO OR3x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR3x2_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.9 1.44 0.972 ; 
        RECT 1.368 0.108 1.44 0.972 ; 
        RECT 1.044 0.108 1.44 0.18 ; 
        RECT 1.044 0.736 1.116 0.972 ; 
        RECT 1.044 0.108 1.116 0.344 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.96 0.972 ; 
      RECT 0.888 0.108 0.96 0.972 ; 
      RECT 0.888 0.504 1.136 0.576 ; 
      RECT 0.16 0.108 0.96 0.18 ; 
  END 
END OR3x2_ASAP7_75t_R 


MACRO OR3x4_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR3x4_ASAP7_75t_R 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.8 ; 
    END 
  END C 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.944 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.9 1.872 0.972 ; 
        RECT 1.8 0.108 1.872 0.972 ; 
        RECT 1.044 0.108 1.872 0.18 ; 
        RECT 1.476 0.736 1.548 0.972 ; 
        RECT 1.476 0.108 1.548 0.344 ; 
        RECT 1.044 0.736 1.116 0.972 ; 
        RECT 1.044 0.108 1.116 0.344 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.16 0.9 0.964 0.972 ; 
      RECT 0.892 0.108 0.964 0.972 ; 
      RECT 0.892 0.504 1.136 0.576 ; 
      RECT 0.16 0.108 0.964 0.18 ; 
  END 
END OR3x4_ASAP7_75t_R 


MACRO OR4x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR4x1_ASAP7_75t_R 0 0 ; 
  SIZE 1.512 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.944 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.944 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.424 0.576 0.944 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.512 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.512 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.272 0.972 ; 
        RECT 0.072 0.108 0.272 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.24 0.9 1.44 0.972 ; 
      RECT 1.368 0.108 1.44 0.972 ; 
      RECT 0.288 0.264 0.36 0.608 ; 
      RECT 0.288 0.264 0.468 0.336 ; 
      RECT 0.396 0.108 0.468 0.336 ; 
      RECT 0.396 0.108 1.44 0.18 ; 
  END 
END OR4x1_ASAP7_75t_R 


MACRO OR4x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR4x2_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.28 1.44 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.28 1.224 0.944 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.944 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.424 0.792 0.944 ; 
    END 
  END D 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.072 0.9 0.488 0.972 ; 
        RECT 0.072 0.108 0.488 0.18 ; 
        RECT 0.072 0.108 0.144 0.972 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 1.456 0.9 1.656 0.972 ; 
      RECT 1.584 0.108 1.656 0.972 ; 
      RECT 0.396 0.252 0.468 0.596 ; 
      RECT 0.396 0.252 0.684 0.324 ; 
      RECT 0.612 0.108 0.684 0.324 ; 
      RECT 0.612 0.108 1.656 0.18 ; 
  END 
END OR4x2_ASAP7_75t_R 


MACRO OR5x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR5x1_ASAP7_75t_R 0 0 ; 
  SIZE 1.728 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.944 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.944 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.944 ; 
    END 
  END D 
  PIN E 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.944 ; 
    END 
  END E 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.728 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.728 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.4 0.9 1.656 0.972 ; 
        RECT 1.584 0.108 1.656 0.972 ; 
        RECT 1.396 0.108 1.656 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.072 0.9 0.28 0.972 ; 
      RECT 0.072 0.108 0.144 0.972 ; 
      RECT 1.368 0.252 1.44 0.616 ; 
      RECT 1.152 0.252 1.44 0.324 ; 
      RECT 1.152 0.108 1.224 0.324 ; 
      RECT 0.072 0.108 1.224 0.18 ; 
  END 
END OR5x1_ASAP7_75t_R 


MACRO OR5x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN OR5x2_ASAP7_75t_R 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.28 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.944 ; 
    END 
  END B 
  PIN C 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.72 0.28 0.792 0.944 ; 
    END 
  END C 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.936 0.28 1.008 0.944 ; 
    END 
  END D 
  PIN E 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.152 0.424 1.224 0.944 ; 
    END 
  END E 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.944 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.456 0.9 1.872 0.972 ; 
        RECT 1.8 0.108 1.872 0.972 ; 
        RECT 1.372 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.072 0.9 0.28 0.972 ; 
      RECT 0.072 0.108 0.144 0.972 ; 
      RECT 1.368 0.252 1.44 0.616 ; 
      RECT 1.152 0.252 1.44 0.324 ; 
      RECT 1.152 0.108 1.224 0.324 ; 
      RECT 0.072 0.108 1.224 0.18 ; 
  END 
END OR5x2_ASAP7_75t_R 


MACRO SDFHx1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFHx1_ASAP7_75t_R 0 0 ; 
  SIZE 5.4 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.396 0.74 0.468 0.944 ; 
        RECT 0.288 0.324 0.468 0.396 ; 
        RECT 0.396 0.136 0.468 0.396 ; 
        RECT 0.288 0.74 0.468 0.812 ; 
        RECT 0.288 0.324 0.36 0.812 ; 
    END 
  END CLK 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.128 0.9 5.328 0.972 ; 
        RECT 5.256 0.108 5.328 0.972 ; 
        RECT 5.128 0.108 5.328 0.18 ; 
    END 
  END QN 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 5.4 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.4 0.036 ; 
    END 
  END VSS 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 1.136 0.432 1.744 0.504 ; 
      LAYER M1 ; 
        RECT 1.584 0.424 1.656 0.656 ; 
      LAYER V1 ; 
        RECT 1.584 0.432 1.656 0.504 ; 
    END 
  END D 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.844 0.144 4.916 0.216 ; 
      LAYER M1 ; 
        RECT 4.824 0.108 5 0.18 ; 
        RECT 4.824 0.108 4.896 0.8 ; 
        RECT 0.864 0.504 1.244 0.576 ; 
        RECT 0.864 0.108 1.032 0.18 ; 
        RECT 0.864 0.108 0.936 0.576 ; 
      LAYER V1 ; 
        RECT 0.864 0.144 0.936 0.216 ; 
        RECT 4.824 0.144 4.896 0.216 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 1.868 0.432 2.36 0.504 ; 
      LAYER M1 ; 
        RECT 1.94 0.756 2.088 0.828 ; 
        RECT 2.016 0.424 2.088 0.828 ; 
        RECT 1.844 0.504 2.088 0.576 ; 
      LAYER V1 ; 
        RECT 2.016 0.432 2.088 0.504 ; 
    END 
  END SI 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.9 4.808 0.972 ; 
      RECT 4.608 0.136 4.68 0.972 ; 
      RECT 4.264 0.9 4.464 0.972 ; 
      RECT 4.392 0.108 4.464 0.972 ; 
      RECT 3.96 0.108 4.032 0.476 ; 
      RECT 3.96 0.108 4.464 0.18 ; 
      RECT 3.616 0.9 3.816 0.972 ; 
      RECT 3.744 0.108 3.816 0.972 ; 
      RECT 3.744 0.612 4.248 0.684 ; 
      RECT 4.176 0.468 4.248 0.684 ; 
      RECT 3.4 0.108 3.816 0.18 ; 
      RECT 3.168 0.9 3.384 0.972 ; 
      RECT 3.312 0.324 3.384 0.972 ; 
      RECT 2.88 0.324 3.384 0.396 ; 
      RECT 3.204 0.18 3.276 0.396 ; 
      RECT 2.88 0.248 2.952 0.396 ; 
      RECT 2.32 0.9 2.808 0.972 ; 
      RECT 2.736 0.108 2.808 0.972 ; 
      RECT 2.736 0.488 3.188 0.56 ; 
      RECT 2.536 0.108 2.808 0.18 ; 
      RECT 2.448 0.612 2.596 0.684 ; 
      RECT 2.448 0.424 2.52 0.684 ; 
      RECT 2.232 0.756 2.38 0.828 ; 
      RECT 2.232 0.424 2.304 0.828 ; 
      RECT 1.044 0.324 1.224 0.396 ; 
      RECT 1.152 0.108 1.224 0.396 ; 
      RECT 1.152 0.108 2 0.18 ; 
      RECT 1.368 0.252 1.44 0.656 ; 
      RECT 1.368 0.252 1.516 0.324 ; 
      RECT 0.592 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.592 0.108 0.792 0.18 ; 
      RECT 0.072 0.9 0.272 0.972 ; 
      RECT 0.072 0.108 0.144 0.972 ; 
      RECT 0.072 0.108 0.272 0.18 ; 
      RECT 5.04 0.36 5.112 0.8 ; 
      RECT 3.528 0.404 3.6 0.668 ; 
      RECT 2.88 0.66 2.952 0.828 ; 
      RECT 1.672 0.252 2.436 0.324 ; 
      RECT 1.02 0.9 2 0.972 ; 
      RECT 1.236 0.756 1.788 0.828 ; 
      RECT 0.504 0.484 0.576 0.668 ; 
    LAYER M2 ; 
      RECT 3.744 0.576 5.132 0.648 ; 
      RECT 1.348 0.288 4.7 0.36 ; 
      RECT 0.052 0.576 3.6 0.648 ; 
      RECT 0.7 0.72 2.972 0.792 ; 
    LAYER V1 ; 
      RECT 5.04 0.576 5.112 0.648 ; 
      RECT 4.608 0.288 4.68 0.36 ; 
      RECT 3.744 0.576 3.816 0.648 ; 
      RECT 3.528 0.576 3.6 0.648 ; 
      RECT 2.88 0.72 2.952 0.792 ; 
      RECT 2.448 0.576 2.52 0.648 ; 
      RECT 2.232 0.72 2.304 0.792 ; 
      RECT 1.368 0.288 1.44 0.36 ; 
      RECT 0.72 0.72 0.792 0.792 ; 
      RECT 0.504 0.576 0.576 0.648 ; 
      RECT 0.072 0.576 0.144 0.648 ; 
  END 
END SDFHx1_ASAP7_75t_R 


MACRO SDFHx2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFHx2_ASAP7_75t_R 0 0 ; 
  SIZE 5.616 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.324 0.468 0.396 ; 
        RECT 0.396 0.136 0.468 0.396 ; 
        RECT 0.288 0.324 0.36 0.8 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.396 1.732 0.468 ; 
        RECT 1.584 0.396 1.656 0.656 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.128 0.9 5.544 0.972 ; 
        RECT 5.472 0.108 5.544 0.972 ; 
        RECT 5.128 0.108 5.544 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.844 0.144 4.916 0.216 ; 
      LAYER M1 ; 
        RECT 4.824 0.108 5 0.18 ; 
        RECT 4.824 0.108 4.896 0.8 ; 
        RECT 0.864 0.504 1.244 0.576 ; 
        RECT 0.864 0.108 1.032 0.18 ; 
        RECT 0.864 0.108 0.936 0.576 ; 
      LAYER V1 ; 
        RECT 0.864 0.144 0.936 0.216 ; 
        RECT 4.824 0.144 4.896 0.216 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.94 0.756 2.088 0.828 ; 
        RECT 2.016 0.424 2.088 0.828 ; 
        RECT 1.844 0.504 2.088 0.576 ; 
    END 
  END SI 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 5.616 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.616 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.9 4.808 0.972 ; 
      RECT 4.608 0.136 4.68 0.972 ; 
      RECT 4.264 0.9 4.464 0.972 ; 
      RECT 4.392 0.108 4.464 0.972 ; 
      RECT 3.96 0.108 4.032 0.476 ; 
      RECT 3.96 0.108 4.464 0.18 ; 
      RECT 3.616 0.9 3.816 0.972 ; 
      RECT 3.744 0.108 3.816 0.972 ; 
      RECT 3.744 0.612 4.248 0.684 ; 
      RECT 4.176 0.468 4.248 0.684 ; 
      RECT 3.4 0.108 3.816 0.18 ; 
      RECT 3.168 0.9 3.384 0.972 ; 
      RECT 3.312 0.324 3.384 0.972 ; 
      RECT 2.88 0.324 3.384 0.396 ; 
      RECT 3.204 0.18 3.276 0.396 ; 
      RECT 2.88 0.248 2.952 0.396 ; 
      RECT 2.32 0.9 2.808 0.972 ; 
      RECT 2.736 0.108 2.808 0.972 ; 
      RECT 2.736 0.488 3.168 0.56 ; 
      RECT 2.536 0.108 2.808 0.18 ; 
      RECT 2.448 0.612 2.596 0.684 ; 
      RECT 2.448 0.424 2.52 0.684 ; 
      RECT 2.232 0.756 2.38 0.828 ; 
      RECT 2.232 0.424 2.304 0.828 ; 
      RECT 1.044 0.324 1.224 0.396 ; 
      RECT 1.152 0.108 1.224 0.396 ; 
      RECT 1.152 0.108 2 0.18 ; 
      RECT 1.368 0.252 1.44 0.656 ; 
      RECT 1.368 0.252 1.516 0.324 ; 
      RECT 0.592 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.592 0.108 0.792 0.18 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.576 0.188 0.648 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 5.04 0.36 5.112 0.8 ; 
      RECT 3.528 0.404 3.6 0.668 ; 
      RECT 2.88 0.66 2.952 0.828 ; 
      RECT 1.672 0.252 2.436 0.324 ; 
      RECT 1.02 0.9 2 0.972 ; 
      RECT 1.236 0.756 1.788 0.828 ; 
      RECT 0.504 0.484 0.576 0.668 ; 
    LAYER M2 ; 
      RECT 3.744 0.576 5.132 0.648 ; 
      RECT 1.348 0.288 4.7 0.36 ; 
      RECT 0.076 0.576 3.6 0.648 ; 
      RECT 0.7 0.72 2.972 0.792 ; 
    LAYER V1 ; 
      RECT 5.04 0.576 5.112 0.648 ; 
      RECT 4.608 0.288 4.68 0.36 ; 
      RECT 3.744 0.576 3.816 0.648 ; 
      RECT 3.528 0.576 3.6 0.648 ; 
      RECT 2.88 0.72 2.952 0.792 ; 
      RECT 2.448 0.576 2.52 0.648 ; 
      RECT 2.232 0.72 2.304 0.792 ; 
      RECT 1.368 0.288 1.44 0.36 ; 
      RECT 0.72 0.72 0.792 0.792 ; 
      RECT 0.504 0.576 0.576 0.648 ; 
      RECT 0.096 0.576 0.168 0.648 ; 
  END 
END SDFHx2_ASAP7_75t_R 


MACRO SDFHx3_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFHx3_ASAP7_75t_R 0 0 ; 
  SIZE 5.832 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.324 0.468 0.396 ; 
        RECT 0.396 0.136 0.468 0.396 ; 
        RECT 0.288 0.324 0.36 0.8 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.396 1.732 0.468 ; 
        RECT 1.584 0.396 1.656 0.656 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.128 0.9 5.76 0.972 ; 
        RECT 5.688 0.108 5.76 0.972 ; 
        RECT 5.128 0.108 5.76 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.844 0.144 4.916 0.216 ; 
      LAYER M1 ; 
        RECT 4.824 0.108 5 0.18 ; 
        RECT 4.824 0.108 4.896 0.8 ; 
        RECT 0.864 0.504 1.244 0.576 ; 
        RECT 0.864 0.108 1.032 0.18 ; 
        RECT 0.864 0.108 0.936 0.576 ; 
      LAYER V1 ; 
        RECT 0.864 0.144 0.936 0.216 ; 
        RECT 4.824 0.144 4.896 0.216 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.94 0.756 2.088 0.828 ; 
        RECT 2.016 0.424 2.088 0.828 ; 
        RECT 1.844 0.504 2.088 0.576 ; 
    END 
  END SI 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 5.832 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.832 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.9 4.808 0.972 ; 
      RECT 4.608 0.136 4.68 0.972 ; 
      RECT 4.264 0.9 4.464 0.972 ; 
      RECT 4.392 0.108 4.464 0.972 ; 
      RECT 3.96 0.108 4.032 0.476 ; 
      RECT 3.96 0.108 4.464 0.18 ; 
      RECT 3.616 0.9 3.816 0.972 ; 
      RECT 3.744 0.108 3.816 0.972 ; 
      RECT 3.744 0.612 4.248 0.684 ; 
      RECT 4.176 0.468 4.248 0.684 ; 
      RECT 3.4 0.108 3.816 0.18 ; 
      RECT 3.168 0.9 3.384 0.972 ; 
      RECT 3.312 0.324 3.384 0.972 ; 
      RECT 2.88 0.324 3.384 0.396 ; 
      RECT 3.204 0.18 3.276 0.396 ; 
      RECT 2.88 0.248 2.952 0.396 ; 
      RECT 2.32 0.9 2.808 0.972 ; 
      RECT 2.736 0.108 2.808 0.972 ; 
      RECT 2.736 0.488 3.168 0.56 ; 
      RECT 2.536 0.108 2.808 0.18 ; 
      RECT 2.448 0.612 2.596 0.684 ; 
      RECT 2.448 0.424 2.52 0.684 ; 
      RECT 2.232 0.756 2.38 0.828 ; 
      RECT 2.232 0.424 2.304 0.828 ; 
      RECT 1.044 0.324 1.224 0.396 ; 
      RECT 1.152 0.108 1.224 0.396 ; 
      RECT 1.152 0.108 2 0.18 ; 
      RECT 1.368 0.252 1.44 0.656 ; 
      RECT 1.368 0.252 1.516 0.324 ; 
      RECT 0.592 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.592 0.108 0.792 0.18 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.576 0.188 0.648 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 5.04 0.36 5.112 0.8 ; 
      RECT 3.528 0.404 3.6 0.668 ; 
      RECT 2.88 0.66 2.952 0.828 ; 
      RECT 1.672 0.252 2.436 0.324 ; 
      RECT 1.02 0.9 2 0.972 ; 
      RECT 1.236 0.756 1.788 0.828 ; 
      RECT 0.504 0.484 0.576 0.668 ; 
    LAYER M2 ; 
      RECT 3.744 0.576 5.132 0.648 ; 
      RECT 1.348 0.288 4.7 0.36 ; 
      RECT 0.076 0.576 3.6 0.648 ; 
      RECT 0.7 0.72 2.972 0.792 ; 
    LAYER V1 ; 
      RECT 5.04 0.576 5.112 0.648 ; 
      RECT 4.608 0.288 4.68 0.36 ; 
      RECT 3.744 0.576 3.816 0.648 ; 
      RECT 3.528 0.576 3.6 0.648 ; 
      RECT 2.88 0.72 2.952 0.792 ; 
      RECT 2.448 0.576 2.52 0.648 ; 
      RECT 2.232 0.72 2.304 0.792 ; 
      RECT 1.368 0.288 1.44 0.36 ; 
      RECT 0.72 0.72 0.792 0.792 ; 
      RECT 0.504 0.576 0.576 0.648 ; 
      RECT 0.096 0.576 0.168 0.648 ; 
  END 
END SDFHx3_ASAP7_75t_R 


MACRO SDFHx4_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFHx4_ASAP7_75t_R 0 0 ; 
  SIZE 6.696 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.252 0.436 0.324 ; 
        RECT 0.288 0.252 0.36 0.8 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.396 1.872 0.656 ; 
        RECT 1.512 0.9 1.836 0.972 ; 
        RECT 1.512 0.396 1.872 0.468 ; 
        RECT 1.512 0.396 1.584 0.972 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.776 0.9 6.624 0.972 ; 
        RECT 6.548 0.108 6.624 0.972 ; 
        RECT 5.776 0.108 6.624 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.916 0.288 2.324 0.36 ; 
      LAYER M1 ; 
        RECT 2.232 0.252 2.396 0.324 ; 
        RECT 2.232 0.252 2.304 0.656 ; 
        RECT 0.936 0.504 1.156 0.576 ; 
        RECT 0.936 0.9 1.084 0.972 ; 
        RECT 0.936 0.108 1.084 0.18 ; 
        RECT 0.936 0.108 1.008 0.972 ; 
      LAYER V1 ; 
        RECT 0.936 0.288 1.008 0.36 ; 
        RECT 2.232 0.288 2.304 0.36 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.772 0.108 3.068 0.18 ; 
        RECT 2.556 0.252 2.844 0.324 ; 
        RECT 2.772 0.108 2.844 0.324 ; 
        RECT 2.448 0.424 2.628 0.496 ; 
        RECT 2.556 0.252 2.628 0.496 ; 
        RECT 2.448 0.424 2.52 0.656 ; 
    END 
  END SI 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 6.696 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.696 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.236 0.9 5.544 0.972 ; 
      RECT 5.472 0.108 5.544 0.972 ; 
      RECT 5.472 0.504 5.788 0.576 ; 
      RECT 4.968 0.504 5.132 0.576 ; 
      RECT 4.968 0.108 5.04 0.576 ; 
      RECT 4.452 0.108 5.544 0.18 ; 
      RECT 4.824 0.728 5.328 0.8 ; 
      RECT 5.256 0.324 5.328 0.8 ; 
      RECT 4.824 0.424 4.896 0.8 ; 
      RECT 5.148 0.324 5.328 0.396 ; 
      RECT 3.528 0.252 3.6 0.656 ; 
      RECT 3.528 0.252 3.924 0.324 ; 
      RECT 3.204 0.9 3.816 0.972 ; 
      RECT 3.744 0.424 3.816 0.972 ; 
      RECT 3.204 0.756 3.276 0.972 ; 
      RECT 2.952 0.756 3.276 0.828 ; 
      RECT 2.952 0.28 3.024 0.828 ; 
      RECT 1.24 0.9 1.44 0.972 ; 
      RECT 1.368 0.108 1.44 0.972 ; 
      RECT 2.016 0.252 2.088 0.656 ; 
      RECT 1.368 0.252 2.088 0.324 ; 
      RECT 1.24 0.108 1.44 0.18 ; 
      RECT 0.592 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.504 0.108 0.792 0.18 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.576 0.188 0.648 ; 
      RECT 0.036 0.108 0.36 0.18 ; 
      RECT 4.608 0.424 4.68 0.8 ; 
      RECT 4.392 0.28 4.464 0.656 ; 
      RECT 4.176 0.424 4.248 0.8 ; 
      RECT 3.312 0.28 3.384 0.668 ; 
      RECT 3.096 0.28 3.168 0.656 ; 
      RECT 2.32 0.9 3.08 0.972 ; 
      RECT 2.736 0.484 2.808 0.668 ; 
      RECT 1.672 0.108 2.648 0.18 ; 
      RECT 1.692 0.756 2.648 0.828 ; 
      RECT 0.504 0.424 0.576 0.8 ; 
    LAYER M2 ; 
      RECT 0.076 0.576 4.7 0.648 ; 
      RECT 0.7 0.432 4.484 0.504 ; 
    LAYER V1 ; 
      RECT 4.608 0.576 4.68 0.648 ; 
      RECT 4.392 0.432 4.464 0.504 ; 
      RECT 4.176 0.576 4.248 0.648 ; 
      RECT 3.312 0.576 3.384 0.648 ; 
      RECT 3.096 0.432 3.168 0.504 ; 
      RECT 2.736 0.576 2.808 0.648 ; 
      RECT 0.72 0.432 0.792 0.504 ; 
      RECT 0.504 0.576 0.576 0.648 ; 
      RECT 0.096 0.576 0.168 0.648 ; 
  END 
END SDFHx4_ASAP7_75t_R 


MACRO SDFLx1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFLx1_ASAP7_75t_R 0 0 ; 
  SIZE 5.4 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.324 0.468 0.396 ; 
        RECT 0.396 0.136 0.468 0.396 ; 
        RECT 0.288 0.324 0.36 0.656 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.396 1.732 0.468 ; 
        RECT 1.584 0.396 1.656 0.656 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.128 0.9 5.328 0.972 ; 
        RECT 5.256 0.108 5.328 0.972 ; 
        RECT 5.128 0.108 5.328 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.844 0.144 4.916 0.216 ; 
      LAYER M1 ; 
        RECT 4.824 0.108 5 0.18 ; 
        RECT 4.824 0.108 4.896 0.8 ; 
        RECT 0.864 0.504 1.244 0.576 ; 
        RECT 0.864 0.108 1.032 0.18 ; 
        RECT 0.864 0.108 0.936 0.576 ; 
      LAYER V1 ; 
        RECT 0.864 0.144 0.936 0.216 ; 
        RECT 4.824 0.144 4.896 0.216 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.94 0.756 2.088 0.828 ; 
        RECT 2.016 0.424 2.088 0.828 ; 
        RECT 1.844 0.504 2.088 0.576 ; 
    END 
  END SI 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 5.4 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.4 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.9 4.808 0.972 ; 
      RECT 4.608 0.136 4.68 0.972 ; 
      RECT 4.264 0.9 4.464 0.972 ; 
      RECT 4.392 0.108 4.464 0.972 ; 
      RECT 3.96 0.108 4.032 0.476 ; 
      RECT 3.96 0.108 4.464 0.18 ; 
      RECT 3.616 0.9 3.816 0.972 ; 
      RECT 3.744 0.108 3.816 0.972 ; 
      RECT 3.744 0.612 4.248 0.684 ; 
      RECT 4.176 0.468 4.248 0.684 ; 
      RECT 3.4 0.108 3.816 0.18 ; 
      RECT 3.168 0.9 3.384 0.972 ; 
      RECT 3.312 0.324 3.384 0.972 ; 
      RECT 2.88 0.324 3.384 0.396 ; 
      RECT 3.204 0.18 3.276 0.396 ; 
      RECT 2.88 0.248 2.952 0.396 ; 
      RECT 2.32 0.9 2.808 0.972 ; 
      RECT 2.736 0.108 2.808 0.972 ; 
      RECT 2.736 0.488 3.188 0.56 ; 
      RECT 2.536 0.108 2.808 0.18 ; 
      RECT 2.448 0.612 2.596 0.684 ; 
      RECT 2.448 0.424 2.52 0.684 ; 
      RECT 2.232 0.756 2.38 0.828 ; 
      RECT 2.232 0.424 2.304 0.828 ; 
      RECT 1.044 0.324 1.224 0.396 ; 
      RECT 1.152 0.108 1.224 0.396 ; 
      RECT 1.152 0.108 2 0.18 ; 
      RECT 1.368 0.252 1.44 0.656 ; 
      RECT 1.368 0.252 1.516 0.324 ; 
      RECT 0.504 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.592 0.108 0.792 0.18 ; 
      RECT 0.428 0.756 0.576 0.828 ; 
      RECT 0.504 0.484 0.576 0.828 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.72 0.188 0.792 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 5.04 0.36 5.112 0.8 ; 
      RECT 3.528 0.404 3.6 0.668 ; 
      RECT 2.88 0.66 2.952 0.828 ; 
      RECT 1.672 0.252 2.436 0.324 ; 
      RECT 1.02 0.9 2 0.972 ; 
      RECT 1.236 0.756 1.788 0.828 ; 
    LAYER M2 ; 
      RECT 3.744 0.576 5.132 0.648 ; 
      RECT 1.348 0.288 4.7 0.36 ; 
      RECT 0.7 0.576 3.6 0.648 ; 
      RECT 0.076 0.72 2.972 0.792 ; 
    LAYER V1 ; 
      RECT 5.04 0.576 5.112 0.648 ; 
      RECT 4.608 0.288 4.68 0.36 ; 
      RECT 3.744 0.576 3.816 0.648 ; 
      RECT 3.528 0.576 3.6 0.648 ; 
      RECT 2.88 0.72 2.952 0.792 ; 
      RECT 2.448 0.576 2.52 0.648 ; 
      RECT 2.232 0.72 2.304 0.792 ; 
      RECT 1.368 0.288 1.44 0.36 ; 
      RECT 0.72 0.576 0.792 0.648 ; 
      RECT 0.504 0.72 0.576 0.792 ; 
      RECT 0.096 0.72 0.168 0.792 ; 
  END 
END SDFLx1_ASAP7_75t_R 


MACRO SDFLx2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFLx2_ASAP7_75t_R 0 0 ; 
  SIZE 5.616 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.324 0.468 0.396 ; 
        RECT 0.396 0.136 0.468 0.396 ; 
        RECT 0.288 0.324 0.36 0.656 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.396 1.732 0.468 ; 
        RECT 1.584 0.396 1.656 0.656 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.128 0.9 5.544 0.972 ; 
        RECT 5.472 0.108 5.544 0.972 ; 
        RECT 5.128 0.108 5.544 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.844 0.144 4.916 0.216 ; 
      LAYER M1 ; 
        RECT 4.824 0.108 5 0.18 ; 
        RECT 4.824 0.108 4.896 0.8 ; 
        RECT 0.864 0.504 1.244 0.576 ; 
        RECT 0.864 0.108 1.032 0.18 ; 
        RECT 0.864 0.108 0.936 0.576 ; 
      LAYER V1 ; 
        RECT 0.864 0.144 0.936 0.216 ; 
        RECT 4.824 0.144 4.896 0.216 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.94 0.756 2.088 0.828 ; 
        RECT 2.016 0.424 2.088 0.828 ; 
        RECT 1.844 0.504 2.088 0.576 ; 
    END 
  END SI 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 5.616 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.616 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.9 4.808 0.972 ; 
      RECT 4.608 0.136 4.68 0.972 ; 
      RECT 4.264 0.9 4.464 0.972 ; 
      RECT 4.392 0.108 4.464 0.972 ; 
      RECT 3.96 0.108 4.032 0.476 ; 
      RECT 3.96 0.108 4.464 0.18 ; 
      RECT 3.616 0.9 3.816 0.972 ; 
      RECT 3.744 0.108 3.816 0.972 ; 
      RECT 3.744 0.612 4.248 0.684 ; 
      RECT 4.176 0.468 4.248 0.684 ; 
      RECT 3.4 0.108 3.816 0.18 ; 
      RECT 3.168 0.9 3.384 0.972 ; 
      RECT 3.312 0.324 3.384 0.972 ; 
      RECT 2.88 0.324 3.384 0.396 ; 
      RECT 3.204 0.18 3.276 0.396 ; 
      RECT 2.88 0.248 2.952 0.396 ; 
      RECT 2.32 0.9 2.808 0.972 ; 
      RECT 2.736 0.108 2.808 0.972 ; 
      RECT 2.736 0.488 3.168 0.56 ; 
      RECT 2.536 0.108 2.808 0.18 ; 
      RECT 2.448 0.612 2.596 0.684 ; 
      RECT 2.448 0.424 2.52 0.684 ; 
      RECT 2.232 0.756 2.38 0.828 ; 
      RECT 2.232 0.424 2.304 0.828 ; 
      RECT 1.044 0.324 1.224 0.396 ; 
      RECT 1.152 0.108 1.224 0.396 ; 
      RECT 1.152 0.108 2 0.18 ; 
      RECT 1.368 0.252 1.44 0.656 ; 
      RECT 1.368 0.252 1.516 0.324 ; 
      RECT 0.504 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.592 0.108 0.792 0.18 ; 
      RECT 0.428 0.756 0.576 0.828 ; 
      RECT 0.504 0.484 0.576 0.828 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.72 0.188 0.792 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 5.04 0.36 5.112 0.8 ; 
      RECT 3.528 0.404 3.6 0.668 ; 
      RECT 2.88 0.66 2.952 0.828 ; 
      RECT 1.672 0.252 2.436 0.324 ; 
      RECT 1.02 0.9 2 0.972 ; 
      RECT 1.236 0.756 1.788 0.828 ; 
    LAYER M2 ; 
      RECT 3.744 0.576 5.132 0.648 ; 
      RECT 1.348 0.288 4.7 0.36 ; 
      RECT 0.7 0.576 3.6 0.648 ; 
      RECT 0.076 0.72 2.972 0.792 ; 
    LAYER V1 ; 
      RECT 5.04 0.576 5.112 0.648 ; 
      RECT 4.608 0.288 4.68 0.36 ; 
      RECT 3.744 0.576 3.816 0.648 ; 
      RECT 3.528 0.576 3.6 0.648 ; 
      RECT 2.88 0.72 2.952 0.792 ; 
      RECT 2.448 0.576 2.52 0.648 ; 
      RECT 2.232 0.72 2.304 0.792 ; 
      RECT 1.368 0.288 1.44 0.36 ; 
      RECT 0.72 0.576 0.792 0.648 ; 
      RECT 0.504 0.72 0.576 0.792 ; 
      RECT 0.096 0.72 0.168 0.792 ; 
  END 
END SDFLx2_ASAP7_75t_R 


MACRO SDFLx3_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFLx3_ASAP7_75t_R 0 0 ; 
  SIZE 5.832 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.324 0.468 0.396 ; 
        RECT 0.396 0.136 0.468 0.396 ; 
        RECT 0.288 0.324 0.36 0.656 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.584 0.396 1.732 0.468 ; 
        RECT 1.584 0.396 1.656 0.656 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.128 0.9 5.76 0.972 ; 
        RECT 5.688 0.108 5.76 0.972 ; 
        RECT 5.128 0.108 5.76 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.844 0.144 4.916 0.216 ; 
      LAYER M1 ; 
        RECT 4.824 0.108 5 0.18 ; 
        RECT 4.824 0.108 4.896 0.8 ; 
        RECT 0.864 0.504 1.244 0.576 ; 
        RECT 0.864 0.108 1.032 0.18 ; 
        RECT 0.864 0.108 0.936 0.576 ; 
      LAYER V1 ; 
        RECT 0.864 0.144 0.936 0.216 ; 
        RECT 4.824 0.144 4.896 0.216 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.94 0.756 2.088 0.828 ; 
        RECT 2.016 0.424 2.088 0.828 ; 
        RECT 1.844 0.504 2.088 0.576 ; 
    END 
  END SI 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 5.832 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 5.832 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.608 0.9 4.808 0.972 ; 
      RECT 4.608 0.136 4.68 0.972 ; 
      RECT 4.264 0.9 4.464 0.972 ; 
      RECT 4.392 0.108 4.464 0.972 ; 
      RECT 3.96 0.108 4.032 0.476 ; 
      RECT 3.96 0.108 4.464 0.18 ; 
      RECT 3.616 0.9 3.816 0.972 ; 
      RECT 3.744 0.108 3.816 0.972 ; 
      RECT 3.744 0.612 4.248 0.684 ; 
      RECT 4.176 0.468 4.248 0.684 ; 
      RECT 3.4 0.108 3.816 0.18 ; 
      RECT 3.168 0.9 3.384 0.972 ; 
      RECT 3.312 0.324 3.384 0.972 ; 
      RECT 2.88 0.324 3.384 0.396 ; 
      RECT 3.204 0.18 3.276 0.396 ; 
      RECT 2.88 0.248 2.952 0.396 ; 
      RECT 2.32 0.9 2.808 0.972 ; 
      RECT 2.736 0.108 2.808 0.972 ; 
      RECT 2.736 0.488 3.168 0.56 ; 
      RECT 2.536 0.108 2.808 0.18 ; 
      RECT 2.448 0.612 2.596 0.684 ; 
      RECT 2.448 0.424 2.52 0.684 ; 
      RECT 2.232 0.756 2.38 0.828 ; 
      RECT 2.232 0.424 2.304 0.828 ; 
      RECT 1.044 0.324 1.224 0.396 ; 
      RECT 1.152 0.108 1.224 0.396 ; 
      RECT 1.152 0.108 2 0.18 ; 
      RECT 1.368 0.252 1.44 0.656 ; 
      RECT 1.368 0.252 1.516 0.324 ; 
      RECT 0.504 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.592 0.108 0.792 0.18 ; 
      RECT 0.428 0.756 0.576 0.828 ; 
      RECT 0.504 0.484 0.576 0.828 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.72 0.188 0.792 ; 
      RECT 0.036 0.108 0.272 0.18 ; 
      RECT 5.04 0.36 5.112 0.8 ; 
      RECT 3.528 0.404 3.6 0.668 ; 
      RECT 2.88 0.66 2.952 0.828 ; 
      RECT 1.672 0.252 2.436 0.324 ; 
      RECT 1.02 0.9 2 0.972 ; 
      RECT 1.236 0.756 1.788 0.828 ; 
    LAYER M2 ; 
      RECT 3.744 0.576 5.132 0.648 ; 
      RECT 1.348 0.288 4.7 0.36 ; 
      RECT 0.7 0.576 3.6 0.648 ; 
      RECT 0.076 0.72 2.972 0.792 ; 
    LAYER V1 ; 
      RECT 5.04 0.576 5.112 0.648 ; 
      RECT 4.608 0.288 4.68 0.36 ; 
      RECT 3.744 0.576 3.816 0.648 ; 
      RECT 3.528 0.576 3.6 0.648 ; 
      RECT 2.88 0.72 2.952 0.792 ; 
      RECT 2.448 0.576 2.52 0.648 ; 
      RECT 2.232 0.72 2.304 0.792 ; 
      RECT 1.368 0.288 1.44 0.36 ; 
      RECT 0.72 0.576 0.792 0.648 ; 
      RECT 0.504 0.72 0.576 0.792 ; 
      RECT 0.096 0.72 0.168 0.792 ; 
  END 
END SDFLx3_ASAP7_75t_R 


MACRO SDFLx4_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN SDFLx4_ASAP7_75t_R 0 0 ; 
  SIZE 6.696 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN CLK 
    DIRECTION INPUT ; 
    USE CLOCK ; 
    PORT 
      LAYER M1 ; 
        RECT 0.288 0.252 0.436 0.324 ; 
        RECT 0.288 0.252 0.36 0.8 ; 
    END 
  END CLK 
  PIN D 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.8 0.396 1.872 0.656 ; 
        RECT 1.512 0.9 1.836 0.972 ; 
        RECT 1.512 0.396 1.872 0.468 ; 
        RECT 1.512 0.396 1.584 0.972 ; 
    END 
  END D 
  PIN QN 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 5.776 0.9 6.624 0.972 ; 
        RECT 6.548 0.108 6.624 0.972 ; 
        RECT 5.776 0.108 6.624 0.18 ; 
    END 
  END QN 
  PIN SE 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.916 0.288 2.324 0.36 ; 
      LAYER M1 ; 
        RECT 2.232 0.252 2.396 0.324 ; 
        RECT 2.232 0.252 2.304 0.656 ; 
        RECT 0.936 0.504 1.156 0.576 ; 
        RECT 0.936 0.9 1.084 0.972 ; 
        RECT 0.936 0.108 1.084 0.18 ; 
        RECT 0.936 0.108 1.008 0.972 ; 
      LAYER V1 ; 
        RECT 0.936 0.288 1.008 0.36 ; 
        RECT 2.232 0.288 2.304 0.36 ; 
    END 
  END SE 
  PIN SI 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 2.772 0.108 3.068 0.18 ; 
        RECT 2.556 0.252 2.844 0.324 ; 
        RECT 2.772 0.108 2.844 0.324 ; 
        RECT 2.448 0.424 2.628 0.496 ; 
        RECT 2.556 0.252 2.628 0.496 ; 
        RECT 2.448 0.424 2.52 0.656 ; 
    END 
  END SI 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 6.696 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 6.696 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 4.236 0.9 5.544 0.972 ; 
      RECT 5.472 0.108 5.544 0.972 ; 
      RECT 5.472 0.504 5.788 0.576 ; 
      RECT 4.968 0.504 5.132 0.576 ; 
      RECT 4.968 0.108 5.04 0.576 ; 
      RECT 4.452 0.108 5.544 0.18 ; 
      RECT 4.824 0.728 5.328 0.8 ; 
      RECT 5.256 0.324 5.328 0.8 ; 
      RECT 4.824 0.424 4.896 0.8 ; 
      RECT 5.148 0.324 5.328 0.396 ; 
      RECT 3.528 0.252 3.6 0.656 ; 
      RECT 3.528 0.252 3.924 0.324 ; 
      RECT 3.204 0.9 3.816 0.972 ; 
      RECT 3.744 0.424 3.816 0.972 ; 
      RECT 3.204 0.756 3.276 0.972 ; 
      RECT 2.952 0.756 3.276 0.828 ; 
      RECT 2.952 0.28 3.024 0.828 ; 
      RECT 1.24 0.9 1.44 0.972 ; 
      RECT 1.368 0.108 1.44 0.972 ; 
      RECT 2.016 0.252 2.088 0.656 ; 
      RECT 1.368 0.252 2.088 0.324 ; 
      RECT 1.24 0.108 1.44 0.18 ; 
      RECT 0.592 0.9 0.792 0.972 ; 
      RECT 0.72 0.108 0.792 0.972 ; 
      RECT 0.504 0.108 0.792 0.18 ; 
      RECT 0.036 0.9 0.272 0.972 ; 
      RECT 0.036 0.108 0.108 0.972 ; 
      RECT 0.036 0.432 0.188 0.504 ; 
      RECT 0.036 0.108 0.36 0.18 ; 
      RECT 4.608 0.424 4.68 0.8 ; 
      RECT 4.392 0.28 4.464 0.656 ; 
      RECT 4.176 0.424 4.248 0.8 ; 
      RECT 3.312 0.28 3.384 0.668 ; 
      RECT 3.096 0.28 3.168 0.656 ; 
      RECT 2.32 0.9 3.08 0.972 ; 
      RECT 2.736 0.484 2.808 0.668 ; 
      RECT 1.672 0.108 2.648 0.18 ; 
      RECT 1.692 0.756 2.648 0.828 ; 
      RECT 0.504 0.412 0.576 0.8 ; 
    LAYER M2 ; 
      RECT 0.7 0.576 4.7 0.648 ; 
      RECT 0.076 0.432 4.484 0.504 ; 
    LAYER V1 ; 
      RECT 4.608 0.576 4.68 0.648 ; 
      RECT 4.392 0.432 4.464 0.504 ; 
      RECT 4.176 0.576 4.248 0.648 ; 
      RECT 3.312 0.576 3.384 0.648 ; 
      RECT 3.096 0.432 3.168 0.504 ; 
      RECT 2.736 0.576 2.808 0.648 ; 
      RECT 0.72 0.576 0.792 0.648 ; 
      RECT 0.504 0.432 0.576 0.504 ; 
      RECT 0.096 0.432 0.168 0.504 ; 
  END 
END SDFLx4_ASAP7_75t_R 


MACRO TAPCELL_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TAPCELL_ASAP7_75t_R 0 0 ; 
  SIZE 0.432 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.432 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.432 0.036 ; 
    END 
  END VSS 
END TAPCELL_ASAP7_75t_R 


MACRO TAPCELL_WITH_FILLER_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TAPCELL_WITH_FILLER_ASAP7_75t_R 0 0 ; 
  SIZE 0.648 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.648 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.648 0.036 ; 
    END 
  END VSS 
END TAPCELL_WITH_FILLER_ASAP7_75t_R 


MACRO TIEHIx1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TIEHIx1_ASAP7_75t_R 0 0 ; 
  SIZE 0.648 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN H 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.376 0.9 0.576 0.972 ; 
        RECT 0.504 0.28 0.576 0.972 ; 
        RECT 0.268 0.28 0.576 0.352 ; 
    END 
  END H 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.648 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.648 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 0.072 0.512 0.38 0.584 ; 
      RECT 0.072 0.108 0.144 0.584 ; 
      RECT 0.072 0.108 0.272 0.18 ; 
  END 
END TIEHIx1_ASAP7_75t_R 


MACRO TIELOx1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN TIELOx1_ASAP7_75t_R 0 0 ; 
  SIZE 0.648 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN L 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.268 0.728 0.576 0.8 ; 
        RECT 0.504 0.108 0.576 0.8 ; 
        RECT 0.376 0.108 0.576 0.18 ; 
    END 
  END L 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 0.648 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 0.648 0.036 ; 
    END 
  END VSS 
  OBS 
    LAYER M1 ; 
      RECT 0.072 0.9 0.272 0.972 ; 
      RECT 0.072 0.496 0.144 0.972 ; 
      RECT 0.072 0.496 0.38 0.568 ; 
  END 
END TIELOx1_ASAP7_75t_R 


MACRO XNOR2x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x1_ASAP7_75t_R 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 1.192 0.288 2.108 0.36 ; 
      LAYER M1 ; 
        RECT 2.016 0.28 2.088 0.608 ; 
        RECT 1.22 0.504 1.46 0.576 ; 
        RECT 1.22 0.268 1.292 0.576 ; 
        RECT 0.852 0.268 1.292 0.34 ; 
        RECT 0.852 0.108 0.924 0.34 ; 
        RECT 0.072 0.108 0.924 0.18 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.108 0.144 0.944 ; 
      LAYER V1 ; 
        RECT 1.22 0.288 1.292 0.36 ; 
        RECT 2.016 0.288 2.088 0.36 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.592 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.9 2.448 0.972 ; 
        RECT 1.8 0.308 1.872 0.972 ; 
        RECT 1.672 0.308 1.872 0.38 ; 
    END 
  END Y 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.484 0.72 2.324 0.792 ; 
      LAYER M1 ; 
        RECT 2.104 0.756 2.304 0.828 ; 
        RECT 2.232 0.484 2.304 0.828 ; 
        RECT 0.428 0.756 0.576 0.828 ; 
        RECT 0.504 0.484 0.576 0.828 ; 
      LAYER V1 ; 
        RECT 0.504 0.72 0.576 0.792 ; 
        RECT 2.232 0.72 2.304 0.792 ; 
    END 
  END A 
  OBS 
    LAYER M1 ; 
      RECT 0.368 0.9 0.772 0.972 ; 
      RECT 0.696 0.756 0.772 0.972 ; 
      RECT 0.696 0.756 1.656 0.828 ; 
      RECT 1.584 0.484 1.656 0.828 ; 
      RECT 0.696 0.328 0.768 0.972 ; 
      RECT 1.024 0.108 2.432 0.18 ; 
  END 
END XNOR2x1_ASAP7_75t_R 


MACRO XNOR2x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.044 0.9 1.76 0.972 ; 
        RECT 1.688 0.504 1.76 0.972 ; 
        RECT 1.564 0.504 1.76 0.576 ; 
        RECT 1.044 0.732 1.116 0.972 ; 
        RECT 0.504 0.732 1.116 0.804 ; 
        RECT 0.504 0.48 0.576 0.804 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.756 1.52 0.828 ; 
        RECT 1.368 0.428 1.44 0.828 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.888 0.9 2.304 0.972 ; 
        RECT 2.232 0.108 2.304 0.972 ; 
        RECT 1.888 0.108 2.304 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.072 0.9 0.252 0.972 ; 
      RECT 0.072 0.108 0.144 0.972 ; 
      RECT 1.908 0.252 1.98 0.604 ; 
      RECT 1.692 0.252 1.98 0.324 ; 
      RECT 1.692 0.108 1.764 0.324 ; 
      RECT 0.072 0.108 1.764 0.18 ; 
      RECT 1.208 0.252 1.28 0.78 ; 
      RECT 0.288 0.252 0.36 0.596 ; 
      RECT 0.288 0.252 1.568 0.324 ; 
      RECT 0.396 0.9 0.92 0.972 ; 
  END 
END XNOR2x2_ASAP7_75t_R 


MACRO XNOR2xp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XNOR2xp5_ASAP7_75t_R 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.252 1.44 0.656 ; 
        RECT 0.828 0.252 1.44 0.324 ; 
        RECT 0.828 0.108 0.9 0.324 ; 
        RECT 0.288 0.108 0.9 0.18 ; 
        RECT 0.288 0.108 0.36 0.8 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.504 0.28 0.576 0.8 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.944 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.9 1.872 0.972 ; 
        RECT 1.8 0.108 1.872 0.972 ; 
        RECT 1.692 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.376 0.9 0.72 0.972 ; 
      RECT 0.648 0.3 0.72 0.972 ; 
      RECT 0.648 0.756 1.656 0.828 ; 
      RECT 1.584 0.484 1.656 0.828 ; 
      RECT 1.044 0.108 1.548 0.18 ; 
  END 
END XNOR2xp5_ASAP7_75t_R 


MACRO XOR2x1_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x1_ASAP7_75t_R 0 0 ; 
  SIZE 2.592 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 1.192 0.72 2.108 0.792 ; 
      LAYER M1 ; 
        RECT 2.016 0.472 2.088 0.8 ; 
        RECT 1.22 0.504 1.46 0.576 ; 
        RECT 0.852 0.74 1.292 0.812 ; 
        RECT 1.22 0.504 1.292 0.812 ; 
        RECT 0.072 0.9 0.924 0.972 ; 
        RECT 0.852 0.74 0.924 0.972 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.136 0.144 0.972 ; 
      LAYER V1 ; 
        RECT 1.22 0.72 1.292 0.792 ; 
        RECT 2.016 0.72 2.088 0.792 ; 
    END 
  END A 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.592 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.592 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.024 0.108 2.448 0.18 ; 
        RECT 1.672 0.7 1.872 0.772 ; 
        RECT 1.8 0.108 1.872 0.772 ; 
    END 
  END Y 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M2 ; 
        RECT 0.484 0.288 2.324 0.36 ; 
      LAYER M1 ; 
        RECT 2.232 0.252 2.304 0.596 ; 
        RECT 2.104 0.252 2.304 0.324 ; 
        RECT 0.504 0.252 0.576 0.596 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
      LAYER V1 ; 
        RECT 0.504 0.288 0.576 0.36 ; 
        RECT 2.232 0.288 2.304 0.36 ; 
    END 
  END B 
  OBS 
    LAYER M1 ; 
      RECT 0.696 0.108 0.768 0.752 ; 
      RECT 1.584 0.252 1.656 0.596 ; 
      RECT 0.696 0.252 1.656 0.324 ; 
      RECT 0.696 0.108 0.772 0.324 ; 
      RECT 0.368 0.108 0.772 0.18 ; 
      RECT 1.024 0.9 2.432 0.972 ; 
  END 
END XOR2x1_ASAP7_75t_R 


MACRO XOR2x2_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2x2_ASAP7_75t_R 0 0 ; 
  SIZE 2.376 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.368 0.252 1.52 0.324 ; 
        RECT 1.368 0.252 1.44 0.652 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.688 0.108 1.76 0.652 ; 
        RECT 1.564 0.504 1.76 0.576 ; 
        RECT 1.044 0.108 1.76 0.18 ; 
        RECT 0.504 0.276 1.116 0.348 ; 
        RECT 1.044 0.108 1.116 0.348 ; 
        RECT 0.504 0.276 0.576 0.6 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 2.376 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 2.376 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.888 0.9 2.304 0.972 ; 
        RECT 2.232 0.108 2.304 0.972 ; 
        RECT 1.888 0.108 2.304 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.072 0.9 1.764 0.972 ; 
      RECT 1.692 0.756 1.764 0.972 ; 
      RECT 0.072 0.108 0.144 0.972 ; 
      RECT 1.692 0.756 1.98 0.828 ; 
      RECT 1.908 0.476 1.98 0.828 ; 
      RECT 0.072 0.108 0.252 0.18 ; 
      RECT 0.288 0.756 1.568 0.828 ; 
      RECT 1.208 0.3 1.28 0.828 ; 
      RECT 0.288 0.484 0.36 0.828 ; 
      RECT 0.396 0.108 0.92 0.18 ; 
  END 
END XOR2x2_ASAP7_75t_R 


MACRO XOR2xp5_ASAP7_75t_R 
  CLASS CORE ; 
  ORIGIN 0 0 ; 
  FOREIGN XOR2xp5_ASAP7_75t_R 0 0 ; 
  SIZE 1.944 BY 1.08 ; 
  SYMMETRY X Y ; 
  SITE asap7sc7p5t ; 
  PIN A 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.828 0.756 1.44 0.828 ; 
        RECT 1.368 0.48 1.44 0.828 ; 
        RECT 0.072 0.9 0.9 0.972 ; 
        RECT 0.828 0.756 0.9 0.972 ; 
        RECT 0.072 0.504 0.312 0.576 ; 
        RECT 0.072 0.136 0.144 0.972 ; 
    END 
  END A 
  PIN B 
    DIRECTION INPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 0.424 0.756 0.576 0.828 ; 
        RECT 0.504 0.252 0.576 0.828 ; 
        RECT 0.428 0.252 0.576 0.324 ; 
    END 
  END B 
  PIN VDD 
    DIRECTION INOUT ; 
    USE POWER ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 1.044 1.944 1.116 ; 
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ; 
    USE GROUND ; 
    SHAPE ABUTMENT ; 
    PORT 
      LAYER M1 ; 
        RECT 0 -0.036 1.944 0.036 ; 
    END 
  END VSS 
  PIN Y 
    DIRECTION OUTPUT ; 
    USE SIGNAL ; 
    PORT 
      LAYER M1 ; 
        RECT 1.692 0.9 1.872 0.972 ; 
        RECT 1.8 0.108 1.872 0.972 ; 
        RECT 1.024 0.108 1.872 0.18 ; 
    END 
  END Y 
  OBS 
    LAYER M1 ; 
      RECT 0.648 0.108 0.72 0.78 ; 
      RECT 1.584 0.252 1.656 0.596 ; 
      RECT 0.648 0.252 1.656 0.324 ; 
      RECT 0.376 0.108 0.72 0.18 ; 
      RECT 1.024 0.9 1.548 0.972 ; 
  END 
END XOR2xp5_ASAP7_75t_R 


END LIBRARY 
